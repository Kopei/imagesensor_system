-- Top_UART_v2.vhd