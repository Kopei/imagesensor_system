-- Version: 9.1 9.1.0.18

library ieee;
use ieee.std_logic_1164.all;
library proasic3;
use proasic3.all;

entity WaveGenSingleZ19 is

    port( RE                      : out   std_logic;
          PLL_Test1_0_SysRst_O    : in    std_logic;
          PLL_Test1_0_Sys_66M_Clk : in    std_logic;
          REen                    : in    std_logic
        );

end WaveGenSingleZ19;

architecture DEF_ARCH of WaveGenSingleZ19 is 

  component OR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component DFN1E1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component XA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OAI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component AX1E
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal CycCnt_n11_0_0_a2_0_0, \CycCnt[10]_net_1\, N_55, 
        \CycCnt[11]_net_1\, CycCnt_n11_0_0_a2_0, 
        \PrState_ns_0_0_a2_0_4[4]\, \PrState_ns_0_0_a2_0_2[4]\, 
        \PrState_ns_0_0_a2_0_1[4]\, N_120, \Phase2Cnt[3]_net_1\, 
        \PrState_ns_0_0_a2_2_4[2]\, \PrState[1]_net_1\, 
        \PrState_ns_0_0_0[2]\, \PrState_ns_0_0_a2_1_0[2]\, 
        \PrState_ns_0_0_a2_1_1[2]\, N_52, 
        \PrState_ns_0_0_a2_2[2]\, \PrState_ns_0_0_a2_0[2]\, 
        CycCntlde_0_a2_2, CycCntlde_0_a2_0, \PrState[2]_net_1\, 
        \PrState[0]_net_1\, \PrState[3]_net_1\, 
        \PrState_ns_0_i_0[1]\, \PrState_ns_0_0_a2_2_7[2]\, N_218, 
        \PrState_ns_0_0_a2_2_6[2]\, \CycCnt[6]_net_1\, 
        \CycCnt[5]_net_1\, \PrState_ns_0_0_a2_2_3[2]\, 
        \PrState_ns_0_0_a2_2_5[2]\, \CycCnt[2]_net_1\, 
        \CycCnt[7]_net_1\, \PrState_ns_0_0_a2_2_1[2]\, 
        \CycCnt[8]_net_1\, \CycCnt[3]_net_1\, \CycCnt[4]_net_1\, 
        \PrState_ns_0_i_a2_0_0[1]\, \PrState_ns_0_i_a2_0_1[1]\, 
        \PrState_ns_0_i_a2_0_0_0[1]\, \PrState_ns_i_0_a2_2[0]\, 
        N_21, \Phase2Cnt[0]_net_1\, \Phase2Cnt[1]_net_1\, N_23, 
        N_212, N_34, N_25, \DelayCnt[5]_net_1\, N_38, N_30, 
        \DelayCnt[2]_net_1\, N_211_i_0, \PrState_ns[2]\, N_11, 
        \Phase1Cnt[0]_net_1\, N_214, N_220, N_215, N_221, N_18, 
        N_231, N_223, N_20, N_22, N_224, N_12, N_219, N_10, N_14, 
        N_54, N_210, N_35, \DelayCnt[4]_net_1\, 
        \DelayCnt[6]_net_1\, \CycCnt[9]_net_1\, N_36, N_88_i_i, 
        N_58, \Phase2Cnt[2]_net_1\, DelayCnt_n0, 
        \DelayCnt[0]_net_1\, \DelayCnt[1]_net_1\, N_27, N_44_i, 
        N_29, \DelayCnt[3]_net_1\, N_60, N_28, N_84, 
        \DelayCnt_RNO_0[3]_net_1\, N_59, \DelayCnt_RNO[4]_net_1\, 
        CycCnt_n9, N_56, CycCnt_n10, N_225, N_81, 
        \CycCnt[1]_net_1\, \CycCnt[0]_net_1\, CycCnt_n11, N_19, 
        CycCnte, CycCnt_n0, \PrState_RNO_4[4]\, \PrState_ns[4]\, 
        N_91, \GND\, \VCC\, GND_0, VCC_0 : std_logic;

begin 


    \CycCnt_RNIEUA[6]\ : OR3C
      port map(A => \CycCnt[5]_net_1\, B => N_221, C => 
        \CycCnt[6]_net_1\, Y => N_223);
    
    WFO : DFN1C0
      port map(D => \PrState[2]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => RE);
    
    \CycCnt[11]\ : DFN1E1C0
      port map(D => CycCnt_n11, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[11]_net_1\);
    
    \PrState[2]\ : DFN1C0
      port map(D => \PrState_ns[2]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \PrState[2]_net_1\);
    
    \PrState_RNO_3[2]\ : NOR2B
      port map(A => \Phase2Cnt[3]_net_1\, B => \PrState[1]_net_1\, 
        Y => \PrState_ns_0_0_a2_0[2]\);
    
    \CycCnt_RNI5Q7[4]\ : NOR2B
      port map(A => N_220, B => \CycCnt[4]_net_1\, Y => N_221);
    
    \DelayCnt[6]\ : DFN1C0
      port map(D => N_27, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \DelayCnt[6]_net_1\);
    
    \DelayCnt_RNI2CRS[1]\ : OR2B
      port map(A => N_212, B => N_36, Y => 
        \PrState_ns_0_i_a2_0_1[1]\);
    
    \CycCnt_RNO_0[6]\ : AO1
      port map(A => N_221, B => \CycCnt[5]_net_1\, C => 
        \CycCnt[6]_net_1\, Y => N_231);
    
    \CycCnt[9]\ : DFN1E1C0
      port map(D => CycCnt_n9, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[9]_net_1\);
    
    \CycCnt_RNO_0[11]\ : OR3A
      port map(A => \CycCnt[10]_net_1\, B => N_55, C => 
        \CycCnt[11]_net_1\, Y => CycCnt_n11_0_0_a2_0_0);
    
    \CycCnt_RNO[7]\ : XA1C
      port map(A => \CycCnt[7]_net_1\, B => N_223, C => N_55, Y
         => N_20);
    
    \PrState_RNO_0[0]\ : NOR3B
      port map(A => \PrState_ns_0_0_a2_0_2[4]\, B => 
        \PrState_ns_0_0_a2_0_1[4]\, C => N_120, Y => 
        \PrState_ns_0_0_a2_0_4[4]\);
    
    \DelayCnt_RNO_0[3]\ : NOR2B
      port map(A => N_34, B => \DelayCnt[2]_net_1\, Y => N_59);
    
    \Phase2Cnt_RNO[2]\ : XA1
      port map(A => N_58, B => \Phase2Cnt[2]_net_1\, C => 
        \PrState[1]_net_1\, Y => N_88_i_i);
    
    \PrState_RNO_4[2]\ : NOR3C
      port map(A => \CycCnt[6]_net_1\, B => \CycCnt[5]_net_1\, C
         => \PrState_ns_0_0_a2_2_3[2]\, Y => 
        \PrState_ns_0_0_a2_2_6[2]\);
    
    \DelayCnt_RNO[1]\ : NOR3A
      port map(A => \PrState[3]_net_1\, B => N_212, C => N_34, Y
         => N_23);
    
    \Phase2Cnt_RNO[1]\ : XA1
      port map(A => \Phase2Cnt[0]_net_1\, B => 
        \Phase2Cnt[1]_net_1\, C => \PrState[1]_net_1\, Y => N_21);
    
    \CycCnt[8]\ : DFN1E1C0
      port map(D => N_22, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[8]_net_1\);
    
    \CycCnt[5]\ : DFN1E1C0
      port map(D => N_215, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[5]_net_1\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \CycCnt_RNO[4]\ : XA1B
      port map(A => \CycCnt[4]_net_1\, B => N_220, C => N_55, Y
         => N_214);
    
    \CycCnt[0]\ : DFN1E1C0
      port map(D => CycCnt_n0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[0]_net_1\);
    
    \PrState_RNI3BM5[2]\ : NOR3B
      port map(A => \Phase2Cnt[3]_net_1\, B => CycCntlde_0_a2_0, 
        C => \PrState[2]_net_1\, Y => CycCntlde_0_a2_2);
    
    \PrState_RNO_1[3]\ : OAI1
      port map(A => N_55, B => \PrState[3]_net_1\, C => REen, Y
         => \PrState_ns_0_i_0[1]\);
    
    \PrState_RNO_10[2]\ : NOR2B
      port map(A => \CycCnt[8]_net_1\, B => \CycCnt[11]_net_1\, Y
         => \PrState_ns_0_0_a2_2_3[2]\);
    
    \DelayCnt_RNI57241[4]\ : NOR2B
      port map(A => N_60, B => \DelayCnt[4]_net_1\, Y => N_38);
    
    \CycCnt_RNO[9]\ : XA1C
      port map(A => \CycCnt[9]_net_1\, B => N_56, C => N_55, Y
         => CycCnt_n9);
    
    \PrState[1]\ : DFN1C0
      port map(D => N_14, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \PrState[1]_net_1\);
    
    \DelayCnt_RNO[4]\ : XA1
      port map(A => \DelayCnt[4]_net_1\, B => N_60, C => 
        \PrState[3]_net_1\, Y => \DelayCnt_RNO[4]_net_1\);
    
    \CycCnt_RNIO9B5[9]\ : NOR2A
      port map(A => \CycCnt[10]_net_1\, B => \CycCnt[9]_net_1\, Y
         => \PrState_ns_0_0_a2_2_4[2]\);
    
    \DelayCnt_RNICHKL[6]\ : OR3B
      port map(A => \DelayCnt[4]_net_1\, B => \DelayCnt[6]_net_1\, 
        C => \DelayCnt[5]_net_1\, Y => \PrState_ns_0_i_a2_0_0[1]\);
    
    \Phase2Cnt_RNIARQC[1]\ : OR3
      port map(A => \Phase2Cnt[0]_net_1\, B => 
        \Phase2Cnt[1]_net_1\, C => \Phase2Cnt[2]_net_1\, Y => 
        N_120);
    
    \DelayCnt_RNIVLDE[1]\ : NOR2B
      port map(A => \DelayCnt[1]_net_1\, B => \DelayCnt[0]_net_1\, 
        Y => N_34);
    
    \CycCnt_RNO[6]\ : NOR3B
      port map(A => N_231, B => N_223, C => N_55, Y => N_18);
    
    \PrState_RNO_0[2]\ : NOR3B
      port map(A => \PrState_ns_0_0_a2_0[2]\, B => REen, C => 
        N_120, Y => \PrState_ns_0_0_a2_2[2]\);
    
    \Phase2Cnt[3]\ : DFN1C0
      port map(D => N_28, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase2Cnt[3]_net_1\);
    
    \PrState_RNIBH0J[4]\ : AO1A
      port map(A => N_120, B => CycCntlde_0_a2_2, C => N_55, Y
         => CycCnte);
    
    \CycCnt_RNIV33[1]\ : NOR2B
      port map(A => \CycCnt[1]_net_1\, B => \CycCnt[0]_net_1\, Y
         => N_218);
    
    \CycCnt[2]\ : DFN1E1C0
      port map(D => N_10, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[2]_net_1\);
    
    \CycCnt_RNO[3]\ : XA1B
      port map(A => \CycCnt[3]_net_1\, B => N_219, C => N_55, Y
         => N_12);
    
    \CycCnt_RNO[2]\ : XA1B
      port map(A => \CycCnt[2]_net_1\, B => N_218, C => N_55, Y
         => N_10);
    
    \PrState_RNO[2]\ : AO1B
      port map(A => \PrState_ns_0_0_a2_2[2]\, B => N_211_i_0, C
         => \PrState_ns_0_0_0[2]\, Y => \PrState_ns[2]\);
    
    \CycCnt_RNO[0]\ : NOR2
      port map(A => N_55, B => \CycCnt[0]_net_1\, Y => CycCnt_n0);
    
    \DelayCnt[2]\ : DFN1C0
      port map(D => N_30, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \DelayCnt[2]_net_1\);
    
    \DelayCnt[5]\ : DFN1C0
      port map(D => N_25, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \DelayCnt[5]_net_1\);
    
    \CycCnt_RNIKGC[7]\ : NOR2A
      port map(A => \CycCnt[7]_net_1\, B => N_223, Y => N_224);
    
    \CycCnt_RNI3LF[9]\ : NOR2A
      port map(A => \CycCnt[9]_net_1\, B => N_56, Y => N_225);
    
    \CycCnt[6]\ : DFN1E1C0
      port map(D => N_18, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[6]_net_1\);
    
    \PrState_RNO_0[1]\ : NOR2
      port map(A => \PrState[1]_net_1\, B => N_35, Y => N_54);
    
    \Phase2Cnt[2]\ : DFN1C0
      port map(D => N_88_i_i, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \Phase2Cnt[2]_net_1\);
    
    \Phase1Cnt[0]\ : DFN1C0
      port map(D => N_35, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[0]_net_1\);
    
    \CycCnt_RNI286[3]\ : NOR2B
      port map(A => N_219, B => \CycCnt[3]_net_1\, Y => N_220);
    
    \DelayCnt[1]\ : DFN1C0
      port map(D => N_23, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \DelayCnt[1]_net_1\);
    
    \PrState_RNIN1U[0]\ : NOR2
      port map(A => \PrState[0]_net_1\, B => \PrState[3]_net_1\, 
        Y => CycCntlde_0_a2_0);
    
    \PrState_RNO_7[2]\ : OR2B
      port map(A => REen, B => \PrState[3]_net_1\, Y => 
        \PrState_ns_0_0_a2_1_0[2]\);
    
    \PrState_RNO_0[3]\ : OR2
      port map(A => N_55, B => \PrState_ns_0_i_a2_0_0[1]\, Y => 
        \PrState_ns_0_i_a2_0_0_0[1]\);
    
    \CycCnt[3]\ : DFN1E1C0
      port map(D => N_12, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[3]_net_1\);
    
    \PrState_RNO_11[2]\ : NOR2B
      port map(A => \CycCnt[3]_net_1\, B => \CycCnt[4]_net_1\, Y
         => \PrState_ns_0_0_a2_2_1[2]\);
    
    \Phase2Cnt_RNO[0]\ : NOR2A
      port map(A => \PrState[1]_net_1\, B => \Phase2Cnt[0]_net_1\, 
        Y => N_29);
    
    \DelayCnt[3]\ : DFN1C0
      port map(D => \DelayCnt_RNO_0[3]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \DelayCnt[3]_net_1\);
    
    \PrState_RNO[1]\ : NOR3A
      port map(A => REen, B => N_54, C => N_210, Y => N_14);
    
    \PrState[4]\ : DFN1P0
      port map(D => \PrState_RNO_4[4]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, PRE => PLL_Test1_0_SysRst_O, Q
         => N_55);
    
    \DelayCnt_RNI2CRS[3]\ : NOR2B
      port map(A => N_36, B => N_34, Y => N_60);
    
    \PrState_RNO_9[2]\ : OR3C
      port map(A => \PrState[2]_net_1\, B => \Phase1Cnt[0]_net_1\, 
        C => REen, Y => N_52);
    
    \Phase2Cnt_RNIROH8[1]\ : NOR2B
      port map(A => \Phase2Cnt[1]_net_1\, B => 
        \Phase2Cnt[0]_net_1\, Y => N_58);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \DelayCnt_RNI3MDE[3]\ : NOR2B
      port map(A => \DelayCnt[3]_net_1\, B => \DelayCnt[2]_net_1\, 
        Y => N_36);
    
    \DelayCnt_RNO[6]\ : NOR2A
      port map(A => \PrState[3]_net_1\, B => N_44_i, Y => N_27);
    
    \CycCnt_RNO[1]\ : XA1B
      port map(A => \CycCnt[0]_net_1\, B => \CycCnt[1]_net_1\, C
         => N_55, Y => N_19);
    
    \CycCnt_RNIR2E[8]\ : OR2B
      port map(A => N_224, B => \CycCnt[8]_net_1\, Y => N_56);
    
    \CycCnt[1]\ : DFN1E1C0
      port map(D => N_19, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[1]_net_1\);
    
    \DelayCnt_RNO[2]\ : XA1
      port map(A => \DelayCnt[2]_net_1\, B => N_34, C => 
        \PrState[3]_net_1\, Y => N_30);
    
    \DelayCnt[4]\ : DFN1C0
      port map(D => \DelayCnt_RNO[4]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \DelayCnt[4]_net_1\);
    
    \CycCnt_RNO[10]\ : XA1B
      port map(A => \CycCnt[10]_net_1\, B => N_225, C => N_55, Y
         => CycCnt_n10);
    
    \DelayCnt_RNO_0[6]\ : AX1E
      port map(A => \DelayCnt[5]_net_1\, B => N_38, C => 
        \DelayCnt[6]_net_1\, Y => N_44_i);
    
    \DelayCnt_RNO[3]\ : XA1
      port map(A => \DelayCnt[3]_net_1\, B => N_59, C => 
        \PrState[3]_net_1\, Y => \DelayCnt_RNO_0[3]_net_1\);
    
    \Phase2Cnt[1]\ : DFN1C0
      port map(D => N_21, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase2Cnt[1]_net_1\);
    
    \PrState_RNO_3[0]\ : NOR2B
      port map(A => \PrState[1]_net_1\, B => REen, Y => 
        \PrState_ns_0_0_a2_0_1[4]\);
    
    \DelayCnt_RNO[5]\ : XA1
      port map(A => \DelayCnt[5]_net_1\, B => N_38, C => 
        \PrState[3]_net_1\, Y => N_25);
    
    \DelayCnt[0]\ : DFN1C0
      port map(D => DelayCnt_n0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \DelayCnt[0]_net_1\);
    
    \CycCnt_RNO_2[11]\ : OR2B
      port map(A => N_225, B => \CycCnt[10]_net_1\, Y => N_81);
    
    \PrState[0]\ : DFN1C0
      port map(D => \PrState_ns[4]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \PrState[0]_net_1\);
    
    \CycCnt_RNO_1[11]\ : NOR2A
      port map(A => \CycCnt[11]_net_1\, B => N_55, Y => 
        CycCnt_n11_0_0_a2_0);
    
    \PrState_RNO_6[2]\ : NOR2B
      port map(A => \PrState_ns_0_0_a2_2_4[2]\, B => N_218, Y => 
        \PrState_ns_0_0_a2_2_7[2]\);
    
    \Phase1Cnt_RNI8TN4[0]\ : NOR2A
      port map(A => \PrState[2]_net_1\, B => \Phase1Cnt[0]_net_1\, 
        Y => N_35);
    
    \PrState_RNO_5[2]\ : NOR3C
      port map(A => \CycCnt[2]_net_1\, B => \CycCnt[7]_net_1\, C
         => \PrState_ns_0_0_a2_2_1[2]\, Y => 
        \PrState_ns_0_0_a2_2_5[2]\);
    
    \CycCnt_RNI0M4[2]\ : NOR2B
      port map(A => N_218, B => \CycCnt[2]_net_1\, Y => N_219);
    
    \CycCnt_RNO[11]\ : MX2A
      port map(A => CycCnt_n11_0_0_a2_0_0, B => 
        CycCnt_n11_0_0_a2_0, S => N_81, Y => CycCnt_n11);
    
    \Phase2Cnt_RNO[3]\ : XA1A
      port map(A => N_84, B => \Phase2Cnt[3]_net_1\, C => 
        \PrState[1]_net_1\, Y => N_28);
    
    \CycCnt[4]\ : DFN1E1C0
      port map(D => N_214, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[4]_net_1\);
    
    \PrState_RNO[3]\ : OA1B
      port map(A => \PrState_ns_0_i_a2_0_1[1]\, B => 
        \PrState_ns_0_i_a2_0_0_0[1]\, C => \PrState_ns_0_i_0[1]\, 
        Y => N_11);
    
    \CycCnt[7]\ : DFN1E1C0
      port map(D => N_20, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[7]_net_1\);
    
    \CycCnt[10]\ : DFN1E1C0
      port map(D => CycCnt_n10, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[10]_net_1\);
    
    \PrState[3]\ : DFN1C0
      port map(D => N_11, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \PrState[3]_net_1\);
    
    \PrState_RNO_1[2]\ : OR3C
      port map(A => \PrState_ns_0_0_a2_2_6[2]\, B => 
        \PrState_ns_0_0_a2_2_5[2]\, C => 
        \PrState_ns_0_0_a2_2_7[2]\, Y => N_211_i_0);
    
    \PrState_RNO[0]\ : AO1A
      port map(A => N_56, B => \PrState_ns_0_0_a2_0_4[4]\, C => 
        N_91, Y => \PrState_ns[4]\);
    
    \Phase2Cnt_RNO_0[3]\ : OR2B
      port map(A => \Phase2Cnt[2]_net_1\, B => N_58, Y => N_84);
    
    \PrState_RNO_0[4]\ : NOR3A
      port map(A => CycCntlde_0_a2_0, B => \PrState[2]_net_1\, C
         => \PrState[1]_net_1\, Y => \PrState_ns_i_0_a2_2[0]\);
    
    \CycCnt_RNO[5]\ : XA1B
      port map(A => \CycCnt[5]_net_1\, B => N_221, C => N_55, Y
         => N_215);
    
    \PrState_RNO_8[2]\ : OR2
      port map(A => \PrState_ns_0_i_a2_0_0[1]\, B => 
        \PrState_ns_0_i_a2_0_1[1]\, Y => 
        \PrState_ns_0_0_a2_1_1[2]\);
    
    \PrState_RNO_2[0]\ : NOR3C
      port map(A => \Phase2Cnt[3]_net_1\, B => \CycCnt[11]_net_1\, 
        C => \PrState_ns_0_0_a2_2_4[2]\, Y => 
        \PrState_ns_0_0_a2_0_2[4]\);
    
    \CycCnt_RNO[8]\ : XA1B
      port map(A => \CycCnt[8]_net_1\, B => N_224, C => N_55, Y
         => N_22);
    
    \PrState_RNO_2[2]\ : OA1
      port map(A => \PrState_ns_0_0_a2_1_0[2]\, B => 
        \PrState_ns_0_0_a2_1_1[2]\, C => N_52, Y => 
        \PrState_ns_0_0_0[2]\);
    
    \PrState_RNO_1[1]\ : NOR3A
      port map(A => \Phase2Cnt[3]_net_1\, B => N_35, C => N_120, 
        Y => N_210);
    
    \Phase2Cnt[0]\ : DFN1C0
      port map(D => N_29, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase2Cnt[0]_net_1\);
    
    \DelayCnt_RNIVLDE_0[1]\ : NOR2
      port map(A => \DelayCnt[1]_net_1\, B => \DelayCnt[0]_net_1\, 
        Y => N_212);
    
    \PrState_RNO[4]\ : OA1C
      port map(A => \PrState_ns_i_0_a2_2[0]\, B => N_55, C => 
        REen, Y => \PrState_RNO_4[4]\);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    \PrState_RNO_1[0]\ : NOR2B
      port map(A => REen, B => \PrState[0]_net_1\, Y => N_91);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    \DelayCnt_RNO[0]\ : NOR2A
      port map(A => \PrState[3]_net_1\, B => \DelayCnt[0]_net_1\, 
        Y => DelayCnt_n0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3;
use proasic3.all;

entity ByteData is

    port( Fifo_dout               : out   std_logic_vector(7 downto 0);
          data_reg_6              : in    std_logic;
          data_reg_0              : in    std_logic;
          data_reg_5              : in    std_logic;
          data_reg_2              : in    std_logic;
          WE                      : in    std_logic;
          RE                      : in    std_logic;
          CMOS_DrvX_0_LVDSen      : in    std_logic;
          ByteData_VCC            : in    std_logic;
          CMOS_DrvX_0_LVDSen_3    : in    std_logic;
          ByteData_GND            : in    std_logic;
          CMOS_DrvX_0_LVDSen_2    : in    std_logic;
          PLL_Test1_0_Sys_66M_Clk : in    std_logic
        );

end ByteData;

architecture DEF_ARCH of ByteData is 

  component AND2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XNOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component RAM4K9
    generic (MEMORYFILE:string := "");

    port( ADDRA11 : in    std_logic := 'U';
          ADDRA10 : in    std_logic := 'U';
          ADDRA9  : in    std_logic := 'U';
          ADDRA8  : in    std_logic := 'U';
          ADDRA7  : in    std_logic := 'U';
          ADDRA6  : in    std_logic := 'U';
          ADDRA5  : in    std_logic := 'U';
          ADDRA4  : in    std_logic := 'U';
          ADDRA3  : in    std_logic := 'U';
          ADDRA2  : in    std_logic := 'U';
          ADDRA1  : in    std_logic := 'U';
          ADDRA0  : in    std_logic := 'U';
          ADDRB11 : in    std_logic := 'U';
          ADDRB10 : in    std_logic := 'U';
          ADDRB9  : in    std_logic := 'U';
          ADDRB8  : in    std_logic := 'U';
          ADDRB7  : in    std_logic := 'U';
          ADDRB6  : in    std_logic := 'U';
          ADDRB5  : in    std_logic := 'U';
          ADDRB4  : in    std_logic := 'U';
          ADDRB3  : in    std_logic := 'U';
          ADDRB2  : in    std_logic := 'U';
          ADDRB1  : in    std_logic := 'U';
          ADDRB0  : in    std_logic := 'U';
          DINA8   : in    std_logic := 'U';
          DINA7   : in    std_logic := 'U';
          DINA6   : in    std_logic := 'U';
          DINA5   : in    std_logic := 'U';
          DINA4   : in    std_logic := 'U';
          DINA3   : in    std_logic := 'U';
          DINA2   : in    std_logic := 'U';
          DINA1   : in    std_logic := 'U';
          DINA0   : in    std_logic := 'U';
          DINB8   : in    std_logic := 'U';
          DINB7   : in    std_logic := 'U';
          DINB6   : in    std_logic := 'U';
          DINB5   : in    std_logic := 'U';
          DINB4   : in    std_logic := 'U';
          DINB3   : in    std_logic := 'U';
          DINB2   : in    std_logic := 'U';
          DINB1   : in    std_logic := 'U';
          DINB0   : in    std_logic := 'U';
          WIDTHA0 : in    std_logic := 'U';
          WIDTHA1 : in    std_logic := 'U';
          WIDTHB0 : in    std_logic := 'U';
          WIDTHB1 : in    std_logic := 'U';
          PIPEA   : in    std_logic := 'U';
          PIPEB   : in    std_logic := 'U';
          WMODEA  : in    std_logic := 'U';
          WMODEB  : in    std_logic := 'U';
          BLKA    : in    std_logic := 'U';
          BLKB    : in    std_logic := 'U';
          WENA    : in    std_logic := 'U';
          WENB    : in    std_logic := 'U';
          CLKA    : in    std_logic := 'U';
          CLKB    : in    std_logic := 'U';
          RESET   : in    std_logic := 'U';
          DOUTA8  : out   std_logic;
          DOUTA7  : out   std_logic;
          DOUTA6  : out   std_logic;
          DOUTA5  : out   std_logic;
          DOUTA4  : out   std_logic;
          DOUTA3  : out   std_logic;
          DOUTA2  : out   std_logic;
          DOUTA1  : out   std_logic;
          DOUTA0  : out   std_logic;
          DOUTB8  : out   std_logic;
          DOUTB7  : out   std_logic;
          DOUTB6  : out   std_logic;
          DOUTB5  : out   std_logic;
          DOUTB4  : out   std_logic;
          DOUTB3  : out   std_logic;
          DOUTB2  : out   std_logic;
          DOUTB1  : out   std_logic;
          DOUTB0  : out   std_logic
        );
  end component;

  component DFN1E1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component INV
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component NAND2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

    signal MEM_RADDR_11_net, RBINNXTSHIFT_11_net, AND2_25_Y, 
        AND2_59_Y, AND2_44_Y, XNOR2_8_Y, MEM_RADDR_7_net, 
        WBINNXTSHIFT_7_net, XOR2_74_Y, MEM_RADDR_12_net, 
        XOR2_36_Y, MEM_RADDR_1_net, MEM_RADDR_9_net, 
        RBINNXTSHIFT_9_net, AO1_21_Y, XOR2_53_Y, AO1_2_Y, 
        AND2_1_Y, RBINNXTSHIFT_2_net, XOR2_34_Y, AO1_14_Y, 
        XNOR2_14_Y, RBINNXTSHIFT_3_net, MEM_WADDR_3_net, 
        XOR2_68_Y, MEM_RADDR_6_net, AO1_4_Y, XOR2_47_Y, AND2_52_Y, 
        AND2_13_Y, NAND2_1_Y, \DFN1P0_EMPTY\, XOR2_0_Y, 
        MEM_WADDR_6_net, AO1_37_Y, XOR2_4_Y, AND2_30_Y, 
        WBINNXTSHIFT_1_net, XOR2_48_Y, AND2_27_Y, AND3_4_Y, 
        XNOR2_15_Y, XNOR2_2_Y, WBINNXTSHIFT_11_net, XOR2_49_Y, 
        AO1_29_Y, MEM_RADDR_10_net, RBINNXTSHIFT_10_net, 
        RAM4K9_QXI_3_DOUTA0, RAM4K9_QXI_3_inst_DOUTA1, 
        RAM4K9_QXI_3_inst_DOUTA2, RAM4K9_QXI_3_inst_DOUTA3, 
        RAM4K9_QXI_3_inst_DOUTA4, RAM4K9_QXI_3_inst_DOUTA5, 
        RAM4K9_QXI_3_inst_DOUTA6, RAM4K9_QXI_3_inst_DOUTA7, 
        RAM4K9_QXI_3_inst_DOUTA8, QXI_3_net, 
        RAM4K9_QXI_3_inst_DOUTB1, RAM4K9_QXI_3_inst_DOUTB2, 
        RAM4K9_QXI_3_inst_DOUTB3, RAM4K9_QXI_3_inst_DOUTB4, 
        RAM4K9_QXI_3_inst_DOUTB5, RAM4K9_QXI_3_inst_DOUTB6, 
        RAM4K9_QXI_3_inst_DOUTB7, RAM4K9_QXI_3_inst_DOUTB8, 
        MEM_WADDR_0_net, MEM_WADDR_1_net, MEM_WADDR_2_net, 
        MEM_WADDR_4_net, MEM_WADDR_5_net, MEM_WADDR_7_net, 
        MEM_WADDR_8_net, MEM_WADDR_9_net, MEM_WADDR_10_net, 
        MEM_WADDR_11_net, MEM_RADDR_0_net, MEM_RADDR_2_net, 
        MEM_RADDR_3_net, MEM_RADDR_4_net, MEM_RADDR_5_net, 
        MEM_RADDR_8_net, MEMWENEG, MEMRENEG, XNOR2_17_Y, AO1_17_Y, 
        XOR2_41_Y, AND2_58_Y, AND2_50_Y, RBINNXTSHIFT_0_net, 
        WBINNXTSHIFT_5_net, AND3_7_Y, XNOR2_12_Y, XNOR2_7_Y, 
        XNOR2_13_Y, AND2_53_Y, XOR2_9_Y, XOR2_3_Y, XOR2_73_Y, 
        RBINNXTSHIFT_1_net, AND2_61_Y, AND2_56_Y, AND2_48_Y, 
        AND2_41_Y, XOR2_66_Y, XOR2_51_Y, AO1_27_Y, XOR2_19_Y, 
        AO1_5_Y, XOR2_76_Y, AO1_36_Y, AND2_8_Y, XNOR2_16_Y, 
        RBINNXTSHIFT_8_net, AO1_25_Y, AO1_23_Y, XNOR2_5_Y, 
        QXI_2_net, DVLDI, XOR2_50_Y, FULLINT, AND3_1_Y, XOR2_40_Y, 
        AND2_4_Y, XOR2_62_Y, XOR2_58_Y, RBINNXTSHIFT_12_net, 
        RAM4K9_QXI_5_DOUTA0, RAM4K9_QXI_5_inst_DOUTA1, 
        RAM4K9_QXI_5_inst_DOUTA2, RAM4K9_QXI_5_inst_DOUTA3, 
        RAM4K9_QXI_5_inst_DOUTA4, RAM4K9_QXI_5_inst_DOUTA5, 
        RAM4K9_QXI_5_inst_DOUTA6, RAM4K9_QXI_5_inst_DOUTA7, 
        RAM4K9_QXI_5_inst_DOUTA8, QXI_5_net, 
        RAM4K9_QXI_5_inst_DOUTB1, RAM4K9_QXI_5_inst_DOUTB2, 
        RAM4K9_QXI_5_inst_DOUTB3, RAM4K9_QXI_5_inst_DOUTB4, 
        RAM4K9_QXI_5_inst_DOUTB5, RAM4K9_QXI_5_inst_DOUTB6, 
        RAM4K9_QXI_5_inst_DOUTB7, RAM4K9_QXI_5_inst_DOUTB8, 
        XOR2_24_Y, AO1_10_Y, AO1_19_Y, AND2_49_Y, AND2_45_Y, 
        XOR2_14_Y, XOR2_65_Y, XOR2_12_Y, MEM_WADDR_12_net, 
        AO1_33_Y, AND2_31_Y, AO1_8_Y, WBINNXTSHIFT_10_net, 
        XOR2_27_Y, AO1_12_Y, XNOR2_23_Y, AO1_16_Y, AND2_26_Y, 
        XOR2_38_Y, WBINNXTSHIFT_6_net, AO1_13_Y, AND2_43_Y, 
        AO1_28_Y, AND2_54_Y, XOR2_16_Y, XOR2_6_Y, XOR2_60_Y, 
        AND2_2_Y, AND2_17_Y, XNOR2_4_Y, AO1_18_Y, AO1_32_Y, 
        XOR2_69_Y, XOR2_7_Y, RBINNXTSHIFT_7_net, XOR2_63_Y, 
        AO1_30_Y, AND2_15_Y, AND2_46_Y, EMPTYINT, XOR2_29_Y, 
        XNOR2_24_Y, RBINNXTSHIFT_4_net, AO1_9_Y, AND2_33_Y, 
        AO1_3_Y, RBINNXTSHIFT_5_net, XOR2_20_Y, AO1_11_Y, 
        AND3_9_Y, XNOR2_18_Y, XNOR2_20_Y, AO1_26_Y, AO1_1_Y, 
        AND2_9_Y, AND2A_0_Y, WBINNXTSHIFT_12_net, AO1_0_Y, 
        AO1_15_Y, AO1_20_Y, AND2_6_Y, MEMORYWE, NAND2_0_Y, 
        XNOR2_10_Y, \DFN1C0_FULL\, AND2_24_Y, AND3_2_Y, AND3_5_Y, 
        AND3_3_Y, AO1_6_Y, XNOR2_22_Y, XOR2_11_Y, XNOR2_3_Y, 
        WBINNXTSHIFT_9_net, RAM4K9_QXI_4_DOUTA0, 
        RAM4K9_QXI_4_inst_DOUTA1, RAM4K9_QXI_4_inst_DOUTA2, 
        RAM4K9_QXI_4_inst_DOUTA3, RAM4K9_QXI_4_inst_DOUTA4, 
        RAM4K9_QXI_4_inst_DOUTA5, RAM4K9_QXI_4_inst_DOUTA6, 
        RAM4K9_QXI_4_inst_DOUTA7, RAM4K9_QXI_4_inst_DOUTA8, 
        QXI_4_net, RAM4K9_QXI_4_inst_DOUTB1, 
        RAM4K9_QXI_4_inst_DOUTB2, RAM4K9_QXI_4_inst_DOUTB3, 
        RAM4K9_QXI_4_inst_DOUTB4, RAM4K9_QXI_4_inst_DOUTB5, 
        RAM4K9_QXI_4_inst_DOUTB6, RAM4K9_QXI_4_inst_DOUTB7, 
        RAM4K9_QXI_4_inst_DOUTB8, WBINNXTSHIFT_3_net, AND2_5_Y, 
        MEMORYRE, WBINNXTSHIFT_2_net, RAM4K9_QXI_0_DOUTA0, 
        RAM4K9_QXI_0_inst_DOUTA1, RAM4K9_QXI_0_inst_DOUTA2, 
        RAM4K9_QXI_0_inst_DOUTA3, RAM4K9_QXI_0_inst_DOUTA4, 
        RAM4K9_QXI_0_inst_DOUTA5, RAM4K9_QXI_0_inst_DOUTA6, 
        RAM4K9_QXI_0_inst_DOUTA7, RAM4K9_QXI_0_inst_DOUTA8, 
        QXI_0_net, RAM4K9_QXI_0_inst_DOUTB1, 
        RAM4K9_QXI_0_inst_DOUTB2, RAM4K9_QXI_0_inst_DOUTB3, 
        RAM4K9_QXI_0_inst_DOUTB4, RAM4K9_QXI_0_inst_DOUTB5, 
        RAM4K9_QXI_0_inst_DOUTB6, RAM4K9_QXI_0_inst_DOUTB7, 
        RAM4K9_QXI_0_inst_DOUTB8, XNOR2_1_Y, WBINNXTSHIFT_0_net, 
        XOR2_10_Y, AO1_24_Y, AND2_3_Y, AND2_10_Y, 
        RBINNXTSHIFT_6_net, XOR2_30_Y, XOR2_22_Y, AND2_19_Y, 
        XOR2_23_Y, AND2_12_Y, AO1_35_Y, XOR2_59_Y, XNOR2_21_Y, 
        RAM4K9_QXI_7_DOUTA0, RAM4K9_QXI_7_inst_DOUTA1, 
        RAM4K9_QXI_7_inst_DOUTA2, RAM4K9_QXI_7_inst_DOUTA3, 
        RAM4K9_QXI_7_inst_DOUTA4, RAM4K9_QXI_7_inst_DOUTA5, 
        RAM4K9_QXI_7_inst_DOUTA6, RAM4K9_QXI_7_inst_DOUTA7, 
        RAM4K9_QXI_7_inst_DOUTA8, QXI_7_net, 
        RAM4K9_QXI_7_inst_DOUTB1, RAM4K9_QXI_7_inst_DOUTB2, 
        RAM4K9_QXI_7_inst_DOUTB3, RAM4K9_QXI_7_inst_DOUTB4, 
        RAM4K9_QXI_7_inst_DOUTB5, RAM4K9_QXI_7_inst_DOUTB6, 
        RAM4K9_QXI_7_inst_DOUTB7, RAM4K9_QXI_7_inst_DOUTB8, 
        XOR2_75_Y, XNOR2_11_Y, AND3_8_Y, AND3_6_Y, AND2_32_Y, 
        AND2_14_Y, XNOR2_6_Y, WBINNXTSHIFT_4_net, AND2_35_Y, 
        QXI_6_net, XOR2_8_Y, WBINNXTSHIFT_8_net, XOR2_72_Y, 
        AO1_34_Y, XNOR2_0_Y, AND2_65_Y, XOR2_1_Y, XNOR2_19_Y, 
        XOR2_61_Y, RAM4K9_QXI_1_DOUTA0, RAM4K9_QXI_1_inst_DOUTA1, 
        RAM4K9_QXI_1_inst_DOUTA2, RAM4K9_QXI_1_inst_DOUTA3, 
        RAM4K9_QXI_1_inst_DOUTA4, RAM4K9_QXI_1_inst_DOUTA5, 
        RAM4K9_QXI_1_inst_DOUTA6, RAM4K9_QXI_1_inst_DOUTA7, 
        RAM4K9_QXI_1_inst_DOUTA8, QXI_1_net, 
        RAM4K9_QXI_1_inst_DOUTB1, RAM4K9_QXI_1_inst_DOUTB2, 
        RAM4K9_QXI_1_inst_DOUTB3, RAM4K9_QXI_1_inst_DOUTB4, 
        RAM4K9_QXI_1_inst_DOUTB5, RAM4K9_QXI_1_inst_DOUTB6, 
        RAM4K9_QXI_1_inst_DOUTB7, RAM4K9_QXI_1_inst_DOUTB8, 
        AND3_0_Y, XNOR2_9_Y, RAM4K9_QXI_2_DOUTA0, 
        RAM4K9_QXI_2_inst_DOUTA1, RAM4K9_QXI_2_inst_DOUTA2, 
        RAM4K9_QXI_2_inst_DOUTA3, RAM4K9_QXI_2_inst_DOUTA4, 
        RAM4K9_QXI_2_inst_DOUTA5, RAM4K9_QXI_2_inst_DOUTA6, 
        RAM4K9_QXI_2_inst_DOUTA7, RAM4K9_QXI_2_inst_DOUTA8, 
        RAM4K9_QXI_2_inst_DOUTB1, RAM4K9_QXI_2_inst_DOUTB2, 
        RAM4K9_QXI_2_inst_DOUTB3, RAM4K9_QXI_2_inst_DOUTB4, 
        RAM4K9_QXI_2_inst_DOUTB5, RAM4K9_QXI_2_inst_DOUTB6, 
        RAM4K9_QXI_2_inst_DOUTB7, RAM4K9_QXI_2_inst_DOUTB8, 
        AO1_7_Y, RAM4K9_QXI_6_DOUTA0, RAM4K9_QXI_6_inst_DOUTA1, 
        RAM4K9_QXI_6_inst_DOUTA2, RAM4K9_QXI_6_inst_DOUTA3, 
        RAM4K9_QXI_6_inst_DOUTA4, RAM4K9_QXI_6_inst_DOUTA5, 
        RAM4K9_QXI_6_inst_DOUTA6, RAM4K9_QXI_6_inst_DOUTA7, 
        RAM4K9_QXI_6_inst_DOUTA8, RAM4K9_QXI_6_inst_DOUTB1, 
        RAM4K9_QXI_6_inst_DOUTB2, RAM4K9_QXI_6_inst_DOUTB3, 
        RAM4K9_QXI_6_inst_DOUTB4, RAM4K9_QXI_6_inst_DOUTB5, 
        RAM4K9_QXI_6_inst_DOUTB6, RAM4K9_QXI_6_inst_DOUTB7, 
        RAM4K9_QXI_6_inst_DOUTB8, \GND\, \VCC\, GND_0, VCC_0
         : std_logic;

begin 


    AND2_2 : AND2
      port map(A => MEM_WADDR_10_net, B => ByteData_GND, Y => 
        AND2_2_Y);
    
    AND3_6 : AND3
      port map(A => XNOR2_14_Y, B => XNOR2_24_Y, C => XNOR2_10_Y, 
        Y => AND3_6_Y);
    
    XNOR2_13 : XNOR2
      port map(A => RBINNXTSHIFT_2_net, B => MEM_WADDR_2_net, Y
         => XNOR2_13_Y);
    
    AO1_11 : AO1
      port map(A => XOR2_10_Y, B => AO1_6_Y, C => AND2_4_Y, Y => 
        AO1_11_Y);
    
    XNOR2_9 : XNOR2
      port map(A => RBINNXTSHIFT_9_net, B => MEM_WADDR_9_net, Y
         => XNOR2_9_Y);
    
    DFN1C0_FULL : DFN1C0
      port map(D => FULLINT, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => CMOS_DrvX_0_LVDSen_2, Q => \DFN1C0_FULL\);
    
    XOR2_19 : XOR2
      port map(A => MEM_WADDR_8_net, B => ByteData_GND, Y => 
        XOR2_19_Y);
    
    AND2_44 : AND2
      port map(A => XOR2_0_Y, B => XOR2_47_Y, Y => AND2_44_Y);
    
    XOR2_23 : XOR2
      port map(A => MEM_RADDR_5_net, B => ByteData_GND, Y => 
        XOR2_23_Y);
    
    XOR2_1 : XOR2
      port map(A => MEM_WADDR_8_net, B => ByteData_GND, Y => 
        XOR2_1_Y);
    
    RAM4K9_QXI_1_inst : RAM4K9
      port map(ADDRA11 => MEM_WADDR_11_net, ADDRA10 => 
        MEM_WADDR_10_net, ADDRA9 => MEM_WADDR_9_net, ADDRA8 => 
        MEM_WADDR_8_net, ADDRA7 => MEM_WADDR_7_net, ADDRA6 => 
        MEM_WADDR_6_net, ADDRA5 => MEM_WADDR_5_net, ADDRA4 => 
        MEM_WADDR_4_net, ADDRA3 => MEM_WADDR_3_net, ADDRA2 => 
        MEM_WADDR_2_net, ADDRA1 => MEM_WADDR_1_net, ADDRA0 => 
        MEM_WADDR_0_net, ADDRB11 => MEM_RADDR_11_net, ADDRB10 => 
        MEM_RADDR_10_net, ADDRB9 => MEM_RADDR_9_net, ADDRB8 => 
        MEM_RADDR_8_net, ADDRB7 => MEM_RADDR_7_net, ADDRB6 => 
        MEM_RADDR_6_net, ADDRB5 => MEM_RADDR_5_net, ADDRB4 => 
        MEM_RADDR_4_net, ADDRB3 => MEM_RADDR_3_net, ADDRB2 => 
        MEM_RADDR_2_net, ADDRB1 => MEM_RADDR_1_net, ADDRB0 => 
        MEM_RADDR_0_net, DINA8 => ByteData_GND, DINA7 => 
        ByteData_GND, DINA6 => ByteData_GND, DINA5 => 
        ByteData_GND, DINA4 => ByteData_GND, DINA3 => 
        ByteData_GND, DINA2 => ByteData_GND, DINA1 => 
        ByteData_GND, DINA0 => ByteData_GND, DINB8 => 
        ByteData_GND, DINB7 => ByteData_GND, DINB6 => 
        ByteData_GND, DINB5 => ByteData_GND, DINB4 => 
        ByteData_GND, DINB3 => ByteData_GND, DINB2 => 
        ByteData_GND, DINB1 => ByteData_GND, DINB0 => 
        ByteData_GND, WIDTHA0 => ByteData_GND, WIDTHA1 => 
        ByteData_GND, WIDTHB0 => ByteData_GND, WIDTHB1 => 
        ByteData_GND, PIPEA => ByteData_GND, PIPEB => 
        ByteData_GND, WMODEA => ByteData_GND, WMODEB => 
        ByteData_GND, BLKA => MEMWENEG, BLKB => MEMRENEG, WENA
         => ByteData_GND, WENB => ByteData_VCC, CLKA => 
        PLL_Test1_0_Sys_66M_Clk, CLKB => PLL_Test1_0_Sys_66M_Clk, 
        RESET => CMOS_DrvX_0_LVDSen, DOUTA8 => 
        RAM4K9_QXI_1_inst_DOUTA8, DOUTA7 => 
        RAM4K9_QXI_1_inst_DOUTA7, DOUTA6 => 
        RAM4K9_QXI_1_inst_DOUTA6, DOUTA5 => 
        RAM4K9_QXI_1_inst_DOUTA5, DOUTA4 => 
        RAM4K9_QXI_1_inst_DOUTA4, DOUTA3 => 
        RAM4K9_QXI_1_inst_DOUTA3, DOUTA2 => 
        RAM4K9_QXI_1_inst_DOUTA2, DOUTA1 => 
        RAM4K9_QXI_1_inst_DOUTA1, DOUTA0 => RAM4K9_QXI_1_DOUTA0, 
        DOUTB8 => RAM4K9_QXI_1_inst_DOUTB8, DOUTB7 => 
        RAM4K9_QXI_1_inst_DOUTB7, DOUTB6 => 
        RAM4K9_QXI_1_inst_DOUTB6, DOUTB5 => 
        RAM4K9_QXI_1_inst_DOUTB5, DOUTB4 => 
        RAM4K9_QXI_1_inst_DOUTB4, DOUTB3 => 
        RAM4K9_QXI_1_inst_DOUTB3, DOUTB2 => 
        RAM4K9_QXI_1_inst_DOUTB2, DOUTB1 => 
        RAM4K9_QXI_1_inst_DOUTB1, DOUTB0 => QXI_1_net);
    
    XOR2_47 : XOR2
      port map(A => MEM_WADDR_7_net, B => ByteData_GND, Y => 
        XOR2_47_Y);
    
    XOR2_38 : XOR2
      port map(A => MEM_WADDR_5_net, B => ByteData_GND, Y => 
        XOR2_38_Y);
    
    AO1_7 : AO1
      port map(A => XOR2_14_Y, B => AO1_18_Y, C => AND2_24_Y, Y
         => AO1_7_Y);
    
    AND2_15 : AND2
      port map(A => MEM_RADDR_2_net, B => ByteData_GND, Y => 
        AND2_15_Y);
    
    AO1_25 : AO1
      port map(A => AND2_54_Y, B => AO1_1_Y, C => AO1_20_Y, Y => 
        AO1_25_Y);
    
    DFN1C0_MEM_WADDR_2_inst : DFN1C0
      port map(D => WBINNXTSHIFT_2_net, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => CMOS_DrvX_0_LVDSen_3, Q
         => MEM_WADDR_2_net);
    
    AND2_1 : AND2
      port map(A => MEM_RADDR_6_net, B => ByteData_GND, Y => 
        AND2_1_Y);
    
    XNOR2_21 : XNOR2
      port map(A => MEM_RADDR_2_net, B => WBINNXTSHIFT_2_net, Y
         => XNOR2_21_Y);
    
    AO1_8 : AO1
      port map(A => XOR2_23_Y, B => AND2_4_Y, C => AND2_14_Y, Y
         => AO1_8_Y);
    
    AND2_49 : AND2
      port map(A => MEM_WADDR_4_net, B => ByteData_GND, Y => 
        AND2_49_Y);
    
    AND2_10 : AND2
      port map(A => MEM_WADDR_5_net, B => ByteData_GND, Y => 
        AND2_10_Y);
    
    XOR2_20 : XOR2
      port map(A => MEM_RADDR_5_net, B => ByteData_GND, Y => 
        XOR2_20_Y);
    
    DFN1E1C0_Q_2_inst : DFN1E1C0
      port map(D => QXI_2_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => CMOS_DrvX_0_LVDSen, E => DVLDI, Q => Fifo_dout(2));
    
    XOR2_63 : XOR2
      port map(A => MEM_RADDR_7_net, B => ByteData_GND, Y => 
        XOR2_63_Y);
    
    XOR2_WBINNXTSHIFT_7_inst : XOR2
      port map(A => XOR2_24_Y, B => AO1_10_Y, Y => 
        WBINNXTSHIFT_7_net);
    
    AND2_12 : AND2
      port map(A => XOR2_60_Y, B => XOR2_22_Y, Y => AND2_12_Y);
    
    AO1_15 : AO1
      port map(A => XOR2_7_Y, B => AND2_26_Y, C => AND2_32_Y, Y
         => AO1_15_Y);
    
    AND2_61 : AND2
      port map(A => MEM_RADDR_0_net, B => MEMORYRE, Y => 
        AND2_61_Y);
    
    AND2_EMPTYINT : AND2
      port map(A => AND3_0_Y, B => XNOR2_22_Y, Y => EMPTYINT);
    
    XOR2_24 : XOR2
      port map(A => MEM_WADDR_7_net, B => ByteData_GND, Y => 
        XOR2_24_Y);
    
    DFN1C0_MEM_WADDR_10_inst : DFN1C0
      port map(D => WBINNXTSHIFT_10_net, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => CMOS_DrvX_0_LVDSen_3, Q
         => MEM_WADDR_10_net);
    
    DFN1C0_MEM_RADDR_0_inst : DFN1C0
      port map(D => RBINNXTSHIFT_0_net, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => CMOS_DrvX_0_LVDSen_2, Q
         => MEM_RADDR_0_net);
    
    DFN1C0_MEM_WADDR_6_inst : DFN1C0
      port map(D => WBINNXTSHIFT_6_net, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => CMOS_DrvX_0_LVDSen_3, Q
         => MEM_WADDR_6_net);
    
    AO1_35 : AO1
      port map(A => XOR2_22_Y, B => AND2_2_Y, C => AND2_5_Y, Y
         => AO1_35_Y);
    
    DFN1E1C0_Q_5_inst : DFN1E1C0
      port map(D => QXI_5_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => CMOS_DrvX_0_LVDSen, E => DVLDI, Q => Fifo_dout(5));
    
    AND2_46 : AND2
      port map(A => MEM_RADDR_3_net, B => ByteData_GND, Y => 
        AND2_46_Y);
    
    XOR2_16 : XOR2
      port map(A => MEM_WADDR_2_net, B => ByteData_GND, Y => 
        XOR2_16_Y);
    
    XOR2_60 : XOR2
      port map(A => MEM_WADDR_10_net, B => ByteData_GND, Y => 
        XOR2_60_Y);
    
    XOR2_RBINNXTSHIFT_7_inst : XOR2
      port map(A => XOR2_63_Y, B => AO1_21_Y, Y => 
        RBINNXTSHIFT_7_net);
    
    AND2_65 : AND2
      port map(A => XNOR2_6_Y, B => XNOR2_11_Y, Y => AND2_65_Y);
    
    AO1_24 : AO1
      port map(A => XOR2_9_Y, B => AO1_14_Y, C => AND2_15_Y, Y
         => AO1_24_Y);
    
    AND2_43 : AND2
      port map(A => AND2_8_Y, B => AND2_12_Y, Y => AND2_43_Y);
    
    AND3_3 : AND3
      port map(A => XNOR2_19_Y, B => XNOR2_0_Y, C => XNOR2_5_Y, Y
         => AND3_3_Y);
    
    RAM4K9_QXI_5_inst : RAM4K9
      port map(ADDRA11 => MEM_WADDR_11_net, ADDRA10 => 
        MEM_WADDR_10_net, ADDRA9 => MEM_WADDR_9_net, ADDRA8 => 
        MEM_WADDR_8_net, ADDRA7 => MEM_WADDR_7_net, ADDRA6 => 
        MEM_WADDR_6_net, ADDRA5 => MEM_WADDR_5_net, ADDRA4 => 
        MEM_WADDR_4_net, ADDRA3 => MEM_WADDR_3_net, ADDRA2 => 
        MEM_WADDR_2_net, ADDRA1 => MEM_WADDR_1_net, ADDRA0 => 
        MEM_WADDR_0_net, ADDRB11 => MEM_RADDR_11_net, ADDRB10 => 
        MEM_RADDR_10_net, ADDRB9 => MEM_RADDR_9_net, ADDRB8 => 
        MEM_RADDR_8_net, ADDRB7 => MEM_RADDR_7_net, ADDRB6 => 
        MEM_RADDR_6_net, ADDRB5 => MEM_RADDR_5_net, ADDRB4 => 
        MEM_RADDR_4_net, ADDRB3 => MEM_RADDR_3_net, ADDRB2 => 
        MEM_RADDR_2_net, ADDRB1 => MEM_RADDR_1_net, ADDRB0 => 
        MEM_RADDR_0_net, DINA8 => ByteData_GND, DINA7 => 
        ByteData_GND, DINA6 => ByteData_GND, DINA5 => 
        ByteData_GND, DINA4 => ByteData_GND, DINA3 => 
        ByteData_GND, DINA2 => ByteData_GND, DINA1 => 
        ByteData_GND, DINA0 => data_reg_5, DINB8 => ByteData_GND, 
        DINB7 => ByteData_GND, DINB6 => ByteData_GND, DINB5 => 
        ByteData_GND, DINB4 => ByteData_GND, DINB3 => 
        ByteData_GND, DINB2 => ByteData_GND, DINB1 => 
        ByteData_GND, DINB0 => ByteData_GND, WIDTHA0 => 
        ByteData_GND, WIDTHA1 => ByteData_GND, WIDTHB0 => 
        ByteData_GND, WIDTHB1 => ByteData_GND, PIPEA => 
        ByteData_GND, PIPEB => ByteData_GND, WMODEA => 
        ByteData_GND, WMODEB => ByteData_GND, BLKA => MEMWENEG, 
        BLKB => MEMRENEG, WENA => ByteData_GND, WENB => 
        ByteData_VCC, CLKA => PLL_Test1_0_Sys_66M_Clk, CLKB => 
        PLL_Test1_0_Sys_66M_Clk, RESET => CMOS_DrvX_0_LVDSen, 
        DOUTA8 => RAM4K9_QXI_5_inst_DOUTA8, DOUTA7 => 
        RAM4K9_QXI_5_inst_DOUTA7, DOUTA6 => 
        RAM4K9_QXI_5_inst_DOUTA6, DOUTA5 => 
        RAM4K9_QXI_5_inst_DOUTA5, DOUTA4 => 
        RAM4K9_QXI_5_inst_DOUTA4, DOUTA3 => 
        RAM4K9_QXI_5_inst_DOUTA3, DOUTA2 => 
        RAM4K9_QXI_5_inst_DOUTA2, DOUTA1 => 
        RAM4K9_QXI_5_inst_DOUTA1, DOUTA0 => RAM4K9_QXI_5_DOUTA0, 
        DOUTB8 => RAM4K9_QXI_5_inst_DOUTB8, DOUTB7 => 
        RAM4K9_QXI_5_inst_DOUTB7, DOUTB6 => 
        RAM4K9_QXI_5_inst_DOUTB6, DOUTB5 => 
        RAM4K9_QXI_5_inst_DOUTB5, DOUTB4 => 
        RAM4K9_QXI_5_inst_DOUTB4, DOUTB3 => 
        RAM4K9_QXI_5_inst_DOUTB3, DOUTB2 => 
        RAM4K9_QXI_5_inst_DOUTB2, DOUTB1 => 
        RAM4K9_QXI_5_inst_DOUTB1, DOUTB0 => QXI_5_net);
    
    MEMWEBUBBLE : INV
      port map(A => MEMORYWE, Y => MEMWENEG);
    
    AND2_6 : AND2
      port map(A => MEM_WADDR_3_net, B => ByteData_GND, Y => 
        AND2_6_Y);
    
    AND3_0 : AND3
      port map(A => XNOR2_9_Y, B => AND3_8_Y, C => AND2_17_Y, Y
         => AND3_0_Y);
    
    XOR2_61 : XOR2
      port map(A => MEM_WADDR_9_net, B => ByteData_GND, Y => 
        XOR2_61_Y);
    
    DFN1E1C0_Q_0_inst : DFN1E1C0
      port map(D => QXI_0_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => CMOS_DrvX_0_LVDSen, E => DVLDI, Q => Fifo_dout(0));
    
    XNOR2_2 : XNOR2
      port map(A => MEM_RADDR_8_net, B => WBINNXTSHIFT_8_net, Y
         => XNOR2_2_Y);
    
    XOR2_49 : XOR2
      port map(A => MEM_WADDR_11_net, B => ByteData_GND, Y => 
        XOR2_49_Y);
    
    XNOR2_19 : XNOR2
      port map(A => MEM_RADDR_3_net, B => WBINNXTSHIFT_3_net, Y
         => XNOR2_19_Y);
    
    AO1_14 : AO1
      port map(A => XOR2_6_Y, B => AND2_61_Y, C => AND2_35_Y, Y
         => AO1_14_Y);
    
    XOR2_WBINNXTSHIFT_2_inst : XOR2
      port map(A => XOR2_11_Y, B => AO1_1_Y, Y => 
        WBINNXTSHIFT_2_net);
    
    XOR2_4 : XOR2
      port map(A => MEM_RADDR_7_net, B => ByteData_GND, Y => 
        XOR2_4_Y);
    
    XOR2_WBINNXTSHIFT_8_inst : XOR2
      port map(A => XOR2_1_Y, B => AO1_5_Y, Y => 
        WBINNXTSHIFT_8_net);
    
    AND3_1 : AND3
      port map(A => XNOR2_3_Y, B => AND3_2_Y, C => AND2_65_Y, Y
         => AND3_1_Y);
    
    AND2_24 : AND2
      port map(A => MEM_RADDR_8_net, B => ByteData_GND, Y => 
        AND2_24_Y);
    
    XOR2_72 : XOR2
      port map(A => MEM_RADDR_4_net, B => ByteData_GND, Y => 
        XOR2_72_Y);
    
    XNOR2_0 : XNOR2
      port map(A => MEM_RADDR_4_net, B => WBINNXTSHIFT_4_net, Y
         => XNOR2_0_Y);
    
    AND2_31 : AND2
      port map(A => XOR2_53_Y, B => XOR2_4_Y, Y => AND2_31_Y);
    
    GND_i : GND
      port map(Y => \GND\);
    
    DFN1C0_MEM_RADDR_12_inst : DFN1C0
      port map(D => RBINNXTSHIFT_12_net, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => CMOS_DrvX_0_LVDSen_2, Q
         => MEM_RADDR_12_net);
    
    XOR2_WBINNXTSHIFT_0_inst : XOR2
      port map(A => MEM_WADDR_0_net, B => MEMORYWE, Y => 
        WBINNXTSHIFT_0_net);
    
    AO1_34 : AO1
      port map(A => AND2_56_Y, B => AO1_18_Y, C => AO1_0_Y, Y => 
        AO1_34_Y);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    DFN1C0_MEM_RADDR_11_inst : DFN1C0
      port map(D => RBINNXTSHIFT_11_net, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => CMOS_DrvX_0_LVDSen_2, Q
         => MEM_RADDR_11_net);
    
    XOR2_8 : XOR2
      port map(A => MEM_RADDR_9_net, B => ByteData_GND, Y => 
        XOR2_8_Y);
    
    XOR2_30 : XOR2
      port map(A => MEM_WADDR_1_net, B => ByteData_GND, Y => 
        XOR2_30_Y);
    
    XOR2_RBINNXTSHIFT_2_inst : XOR2
      port map(A => XOR2_34_Y, B => AO1_14_Y, Y => 
        RBINNXTSHIFT_2_net);
    
    XOR2_RBINNXTSHIFT_8_inst : XOR2
      port map(A => XOR2_73_Y, B => AO1_18_Y, Y => 
        RBINNXTSHIFT_8_net);
    
    MEMREBUBBLE : INV
      port map(A => MEMORYRE, Y => MEMRENEG);
    
    AND2_35 : AND2
      port map(A => MEM_RADDR_1_net, B => ByteData_GND, Y => 
        AND2_35_Y);
    
    XOR2_RBINNXTSHIFT_0_inst : XOR2
      port map(A => MEM_RADDR_0_net, B => MEMORYRE, Y => 
        RBINNXTSHIFT_0_net);
    
    XOR2_34 : XOR2
      port map(A => MEM_RADDR_2_net, B => ByteData_GND, Y => 
        XOR2_34_Y);
    
    XOR2_WBINNXTSHIFT_1_inst : XOR2
      port map(A => XOR2_48_Y, B => AND2_27_Y, Y => 
        WBINNXTSHIFT_1_net);
    
    AND2_3 : AND2
      port map(A => AND2_19_Y, B => AND2_31_Y, Y => AND2_3_Y);
    
    AND2_30 : AND2
      port map(A => MEM_RADDR_7_net, B => ByteData_GND, Y => 
        AND2_30_Y);
    
    XNOR2_6 : XNOR2
      port map(A => MEM_RADDR_10_net, B => WBINNXTSHIFT_10_net, Y
         => XNOR2_6_Y);
    
    AND2_14 : AND2
      port map(A => MEM_RADDR_5_net, B => ByteData_GND, Y => 
        AND2_14_Y);
    
    XOR2_RBINNXTSHIFT_10_inst : XOR2
      port map(A => XOR2_29_Y, B => AO1_16_Y, Y => 
        RBINNXTSHIFT_10_net);
    
    AND2_32 : AND2
      port map(A => MEM_RADDR_11_net, B => ByteData_GND, Y => 
        AND2_32_Y);
    
    AND3_8 : AND3
      port map(A => AND3_9_Y, B => AND3_7_Y, C => AND3_6_Y, Y => 
        AND3_8_Y);
    
    DFN1C0_MEM_WADDR_5_inst : DFN1C0
      port map(D => WBINNXTSHIFT_5_net, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => CMOS_DrvX_0_LVDSen_3, Q
         => MEM_WADDR_5_net);
    
    XNOR2_11 : XNOR2
      port map(A => MEM_RADDR_11_net, B => WBINNXTSHIFT_11_net, Y
         => XNOR2_11_Y);
    
    AO1_2 : AO1
      port map(A => AND2_19_Y, B => AO1_6_Y, C => AO1_8_Y, Y => 
        AO1_2_Y);
    
    XOR2_75 : XOR2
      port map(A => MEM_WADDR_4_net, B => ByteData_GND, Y => 
        XOR2_75_Y);
    
    AND2_26 : AND2
      port map(A => MEM_RADDR_10_net, B => ByteData_GND, Y => 
        AND2_26_Y);
    
    XOR2_9 : XOR2
      port map(A => MEM_RADDR_2_net, B => ByteData_GND, Y => 
        XOR2_9_Y);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    AND3_5 : AND3
      port map(A => XNOR2_1_Y, B => XNOR2_17_Y, C => XNOR2_21_Y, 
        Y => AND3_5_Y);
    
    RAM4K9_QXI_4_inst : RAM4K9
      port map(ADDRA11 => MEM_WADDR_11_net, ADDRA10 => 
        MEM_WADDR_10_net, ADDRA9 => MEM_WADDR_9_net, ADDRA8 => 
        MEM_WADDR_8_net, ADDRA7 => MEM_WADDR_7_net, ADDRA6 => 
        MEM_WADDR_6_net, ADDRA5 => MEM_WADDR_5_net, ADDRA4 => 
        MEM_WADDR_4_net, ADDRA3 => MEM_WADDR_3_net, ADDRA2 => 
        MEM_WADDR_2_net, ADDRA1 => MEM_WADDR_1_net, ADDRA0 => 
        MEM_WADDR_0_net, ADDRB11 => MEM_RADDR_11_net, ADDRB10 => 
        MEM_RADDR_10_net, ADDRB9 => MEM_RADDR_9_net, ADDRB8 => 
        MEM_RADDR_8_net, ADDRB7 => MEM_RADDR_7_net, ADDRB6 => 
        MEM_RADDR_6_net, ADDRB5 => MEM_RADDR_5_net, ADDRB4 => 
        MEM_RADDR_4_net, ADDRB3 => MEM_RADDR_3_net, ADDRB2 => 
        MEM_RADDR_2_net, ADDRB1 => MEM_RADDR_1_net, ADDRB0 => 
        MEM_RADDR_0_net, DINA8 => ByteData_GND, DINA7 => 
        ByteData_GND, DINA6 => ByteData_GND, DINA5 => 
        ByteData_GND, DINA4 => ByteData_GND, DINA3 => 
        ByteData_GND, DINA2 => ByteData_GND, DINA1 => 
        ByteData_GND, DINA0 => ByteData_GND, DINB8 => 
        ByteData_GND, DINB7 => ByteData_GND, DINB6 => 
        ByteData_GND, DINB5 => ByteData_GND, DINB4 => 
        ByteData_GND, DINB3 => ByteData_GND, DINB2 => 
        ByteData_GND, DINB1 => ByteData_GND, DINB0 => 
        ByteData_GND, WIDTHA0 => ByteData_GND, WIDTHA1 => 
        ByteData_GND, WIDTHB0 => ByteData_GND, WIDTHB1 => 
        ByteData_GND, PIPEA => ByteData_GND, PIPEB => 
        ByteData_GND, WMODEA => ByteData_GND, WMODEB => 
        ByteData_GND, BLKA => MEMWENEG, BLKB => MEMRENEG, WENA
         => ByteData_GND, WENB => ByteData_VCC, CLKA => 
        PLL_Test1_0_Sys_66M_Clk, CLKB => PLL_Test1_0_Sys_66M_Clk, 
        RESET => CMOS_DrvX_0_LVDSen, DOUTA8 => 
        RAM4K9_QXI_4_inst_DOUTA8, DOUTA7 => 
        RAM4K9_QXI_4_inst_DOUTA7, DOUTA6 => 
        RAM4K9_QXI_4_inst_DOUTA6, DOUTA5 => 
        RAM4K9_QXI_4_inst_DOUTA5, DOUTA4 => 
        RAM4K9_QXI_4_inst_DOUTA4, DOUTA3 => 
        RAM4K9_QXI_4_inst_DOUTA3, DOUTA2 => 
        RAM4K9_QXI_4_inst_DOUTA2, DOUTA1 => 
        RAM4K9_QXI_4_inst_DOUTA1, DOUTA0 => RAM4K9_QXI_4_DOUTA0, 
        DOUTB8 => RAM4K9_QXI_4_inst_DOUTB8, DOUTB7 => 
        RAM4K9_QXI_4_inst_DOUTB7, DOUTB6 => 
        RAM4K9_QXI_4_inst_DOUTB6, DOUTB5 => 
        RAM4K9_QXI_4_inst_DOUTB5, DOUTB4 => 
        RAM4K9_QXI_4_inst_DOUTB4, DOUTB3 => 
        RAM4K9_QXI_4_inst_DOUTB3, DOUTB2 => 
        RAM4K9_QXI_4_inst_DOUTB2, DOUTB1 => 
        RAM4K9_QXI_4_inst_DOUTB1, DOUTB0 => QXI_4_net);
    
    XOR2_RBINNXTSHIFT_1_inst : XOR2
      port map(A => XOR2_36_Y, B => AND2_61_Y, Y => 
        RBINNXTSHIFT_1_net);
    
    XOR2_59 : XOR2
      port map(A => MEM_WADDR_6_net, B => ByteData_GND, Y => 
        XOR2_59_Y);
    
    XNOR2_4 : XNOR2
      port map(A => RBINNXTSHIFT_11_net, B => MEM_WADDR_11_net, Y
         => XNOR2_4_Y);
    
    XNOR2_20 : XNOR2
      port map(A => RBINNXTSHIFT_7_net, B => MEM_WADDR_7_net, Y
         => XNOR2_20_Y);
    
    DFN1E1C0_Q_1_inst : DFN1E1C0
      port map(D => QXI_1_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => CMOS_DrvX_0_LVDSen, E => DVLDI, Q => Fifo_dout(1));
    
    DFN1C0_MEM_RADDR_7_inst : DFN1C0
      port map(D => RBINNXTSHIFT_7_net, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => CMOS_DrvX_0_LVDSen_3, Q
         => MEM_RADDR_7_net);
    
    DFN1C0_MEM_WADDR_4_inst : DFN1C0
      port map(D => WBINNXTSHIFT_4_net, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => CMOS_DrvX_0_LVDSen_3, Q
         => MEM_WADDR_4_net);
    
    XOR2_WBINNXTSHIFT_10_inst : XOR2
      port map(A => XOR2_27_Y, B => AO1_12_Y, Y => 
        WBINNXTSHIFT_10_net);
    
    AO1_28 : AO1
      port map(A => AND2_12_Y, B => AO1_17_Y, C => AO1_35_Y, Y
         => AO1_28_Y);
    
    AND2_19 : AND2
      port map(A => XOR2_10_Y, B => XOR2_23_Y, Y => AND2_19_Y);
    
    DFN1C0_MEM_WADDR_8_inst : DFN1C0
      port map(D => WBINNXTSHIFT_8_net, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => CMOS_DrvX_0_LVDSen_3, Q
         => MEM_WADDR_8_net);
    
    XOR2_22 : XOR2
      port map(A => MEM_WADDR_11_net, B => ByteData_GND, Y => 
        XOR2_22_Y);
    
    AO1_1 : AO1
      port map(A => XOR2_30_Y, B => AND2_27_Y, C => AND2_45_Y, Y
         => AO1_1_Y);
    
    DFN1E1C0_Q_4_inst : DFN1E1C0
      port map(D => QXI_4_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => CMOS_DrvX_0_LVDSen, E => DVLDI, Q => Fifo_dout(4));
    
    XNOR2_18 : XNOR2
      port map(A => RBINNXTSHIFT_6_net, B => MEM_WADDR_6_net, Y
         => XNOR2_18_Y);
    
    XOR2_WBINNXTSHIFT_3_inst : XOR2
      port map(A => XOR2_69_Y, B => AO1_26_Y, Y => 
        WBINNXTSHIFT_3_net);
    
    AO1_3 : AO1
      port map(A => XOR2_58_Y, B => AND2_49_Y, C => AND2_10_Y, Y
         => AO1_3_Y);
    
    DFN1C0_MEM_RADDR_6_inst : DFN1C0
      port map(D => RBINNXTSHIFT_6_net, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => CMOS_DrvX_0_LVDSen_3, Q
         => MEM_RADDR_6_net);
    
    AO1_18 : AO1
      port map(A => AND2_3_Y, B => AO1_6_Y, C => AO1_33_Y, Y => 
        AO1_18_Y);
    
    XOR2_48 : XOR2
      port map(A => MEM_WADDR_1_net, B => ByteData_GND, Y => 
        XOR2_48_Y);
    
    DFN1E1C0_Q_7_inst : DFN1E1C0
      port map(D => QXI_7_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => CMOS_DrvX_0_LVDSen, E => DVLDI, Q => Fifo_dout(7));
    
    XOR2_62 : XOR2
      port map(A => MEM_WADDR_4_net, B => ByteData_GND, Y => 
        XOR2_62_Y);
    
    AND2_13 : AND2
      port map(A => MEM_WADDR_7_net, B => ByteData_GND, Y => 
        AND2_13_Y);
    
    XOR2_10 : XOR2
      port map(A => MEM_RADDR_4_net, B => ByteData_GND, Y => 
        XOR2_10_Y);
    
    XNOR2_1 : XNOR2
      port map(A => MEM_RADDR_0_net, B => WBINNXTSHIFT_0_net, Y
         => XNOR2_1_Y);
    
    AND2_58 : AND2
      port map(A => MEM_WADDR_8_net, B => ByteData_GND, Y => 
        AND2_58_Y);
    
    XOR2_RBINNXTSHIFT_3_inst : XOR2
      port map(A => XOR2_51_Y, B => AO1_24_Y, Y => 
        RBINNXTSHIFT_3_net);
    
    XOR2_27 : XOR2
      port map(A => MEM_WADDR_10_net, B => ByteData_GND, Y => 
        XOR2_27_Y);
    
    AND2_MEMORYRE : AND2
      port map(A => NAND2_1_Y, B => RE, Y => MEMORYRE);
    
    XOR2_7 : XOR2
      port map(A => MEM_RADDR_11_net, B => ByteData_GND, Y => 
        XOR2_7_Y);
    
    AND2_5 : AND2
      port map(A => MEM_WADDR_11_net, B => ByteData_GND, Y => 
        AND2_5_Y);
    
    XOR2_14 : XOR2
      port map(A => MEM_RADDR_8_net, B => ByteData_GND, Y => 
        XOR2_14_Y);
    
    AND2_50 : AND2
      port map(A => MEM_WADDR_9_net, B => ByteData_GND, Y => 
        AND2_50_Y);
    
    XOR2_11 : XOR2
      port map(A => MEM_WADDR_2_net, B => ByteData_GND, Y => 
        XOR2_11_Y);
    
    XNOR2_3 : XNOR2
      port map(A => MEM_RADDR_9_net, B => WBINNXTSHIFT_9_net, Y
         => XNOR2_3_Y);
    
    XNOR2_22 : XNOR2
      port map(A => RBINNXTSHIFT_12_net, B => MEM_WADDR_12_net, Y
         => XNOR2_22_Y);
    
    AND2_52 : AND2
      port map(A => MEM_WADDR_6_net, B => ByteData_GND, Y => 
        AND2_52_Y);
    
    XNOR2_15 : XNOR2
      port map(A => MEM_RADDR_6_net, B => WBINNXTSHIFT_6_net, Y
         => XNOR2_15_Y);
    
    DFN1C0_MEM_RADDR_3_inst : DFN1C0
      port map(D => RBINNXTSHIFT_3_net, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => CMOS_DrvX_0_LVDSen_3, Q
         => MEM_RADDR_3_net);
    
    XOR2_WBINNXTSHIFT_9_inst : XOR2
      port map(A => XOR2_61_Y, B => AO1_27_Y, Y => 
        WBINNXTSHIFT_9_net);
    
    AO1_6 : AO1
      port map(A => AND2_53_Y, B => AO1_14_Y, C => AO1_30_Y, Y
         => AO1_6_Y);
    
    XOR2_WBINNXTSHIFT_4_inst : XOR2
      port map(A => XOR2_75_Y, B => AO1_25_Y, Y => 
        WBINNXTSHIFT_4_net);
    
    AND3_2 : AND3
      port map(A => AND3_4_Y, B => AND3_5_Y, C => AND3_3_Y, Y => 
        AND3_2_Y);
    
    AO1_12 : AO1
      port map(A => AND2_8_Y, B => AO1_5_Y, C => AO1_17_Y, Y => 
        AO1_12_Y);
    
    AND2_9 : AND2
      port map(A => MEM_WADDR_2_net, B => ByteData_GND, Y => 
        AND2_9_Y);
    
    XOR2_65 : XOR2
      port map(A => MEM_RADDR_9_net, B => ByteData_GND, Y => 
        XOR2_65_Y);
    
    XOR2_58 : XOR2
      port map(A => MEM_WADDR_5_net, B => ByteData_GND, Y => 
        XOR2_58_Y);
    
    DFN1C0_MEM_WADDR_1_inst : DFN1C0
      port map(D => WBINNXTSHIFT_1_net, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => CMOS_DrvX_0_LVDSen_3, Q
         => MEM_WADDR_1_net);
    
    AO1_32 : AO1
      port map(A => XOR2_65_Y, B => AND2_24_Y, C => AND2_33_Y, Y
         => AO1_32_Y);
    
    AO1_9 : AO1
      port map(A => AND2_59_Y, B => AO1_25_Y, C => AO1_3_Y, Y => 
        AO1_9_Y);
    
    XOR2_RBINNXTSHIFT_9_inst : XOR2
      port map(A => XOR2_8_Y, B => AO1_7_Y, Y => 
        RBINNXTSHIFT_9_net);
    
    NAND2_0 : NAND2
      port map(A => \DFN1C0_FULL\, B => ByteData_VCC, Y => 
        NAND2_0_Y);
    
    DFN1C0_MEM_RADDR_10_inst : DFN1C0
      port map(D => RBINNXTSHIFT_10_net, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => CMOS_DrvX_0_LVDSen_2, Q
         => MEM_RADDR_10_net);
    
    DFN1E1C0_Q_3_inst : DFN1E1C0
      port map(D => QXI_3_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => CMOS_DrvX_0_LVDSen, E => DVLDI, Q => Fifo_dout(3));
    
    XOR2_RBINNXTSHIFT_4_inst : XOR2
      port map(A => XOR2_72_Y, B => AO1_6_Y, Y => 
        RBINNXTSHIFT_4_net);
    
    XOR2_76 : XOR2
      port map(A => MEM_RADDR_11_net, B => ByteData_GND, Y => 
        XOR2_76_Y);
    
    AND2_27 : AND2
      port map(A => MEM_WADDR_0_net, B => MEMORYWE, Y => 
        AND2_27_Y);
    
    DFN1C0_MEM_RADDR_5_inst : DFN1C0
      port map(D => RBINNXTSHIFT_5_net, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => CMOS_DrvX_0_LVDSen_3, Q
         => MEM_RADDR_5_net);
    
    DFN1C0_DVLDI : DFN1C0
      port map(D => AND2A_0_Y, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => CMOS_DrvX_0_LVDSen_2, Q => DVLDI);
    
    XNOR2_10 : XNOR2
      port map(A => RBINNXTSHIFT_5_net, B => MEM_WADDR_5_net, Y
         => XNOR2_10_Y);
    
    AO1_20 : AO1
      port map(A => XOR2_66_Y, B => AND2_9_Y, C => AND2_6_Y, Y
         => AO1_20_Y);
    
    AND2_MEMORYWE : AND2
      port map(A => NAND2_0_Y, B => WE, Y => MEMORYWE);
    
    DFN1C0_MEM_WADDR_9_inst : DFN1C0
      port map(D => WBINNXTSHIFT_9_net, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => CMOS_DrvX_0_LVDSen_3, Q
         => MEM_WADDR_9_net);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    AO1_0 : AO1
      port map(A => AND2_41_Y, B => AO1_32_Y, C => AO1_15_Y, Y
         => AO1_0_Y);
    
    XOR2_29 : XOR2
      port map(A => MEM_RADDR_10_net, B => ByteData_GND, Y => 
        XOR2_29_Y);
    
    XOR2_40 : XOR2
      port map(A => MEM_RADDR_12_net, B => WBINNXTSHIFT_12_net, Y
         => XOR2_40_Y);
    
    DFN1C0_MEM_WADDR_0_inst : DFN1C0
      port map(D => WBINNXTSHIFT_0_net, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => CMOS_DrvX_0_LVDSen_3, Q
         => MEM_WADDR_0_net);
    
    AND2A_0 : AND2A
      port map(A => \DFN1P0_EMPTY\, B => RE, Y => AND2A_0_Y);
    
    AO1_26 : AO1
      port map(A => XOR2_16_Y, B => AO1_1_Y, C => AND2_9_Y, Y => 
        AO1_26_Y);
    
    AND3_9 : AND3
      port map(A => XNOR2_18_Y, B => XNOR2_20_Y, C => XNOR2_16_Y, 
        Y => AND3_9_Y);
    
    AO1_23 : AO1
      port map(A => AND2_44_Y, B => AO1_3_Y, C => AO1_4_Y, Y => 
        AO1_23_Y);
    
    AND2_33 : AND2
      port map(A => MEM_RADDR_9_net, B => ByteData_GND, Y => 
        AND2_33_Y);
    
    RAM4K9_QXI_0_inst : RAM4K9
      port map(ADDRA11 => MEM_WADDR_11_net, ADDRA10 => 
        MEM_WADDR_10_net, ADDRA9 => MEM_WADDR_9_net, ADDRA8 => 
        MEM_WADDR_8_net, ADDRA7 => MEM_WADDR_7_net, ADDRA6 => 
        MEM_WADDR_6_net, ADDRA5 => MEM_WADDR_5_net, ADDRA4 => 
        MEM_WADDR_4_net, ADDRA3 => MEM_WADDR_3_net, ADDRA2 => 
        MEM_WADDR_2_net, ADDRA1 => MEM_WADDR_1_net, ADDRA0 => 
        MEM_WADDR_0_net, ADDRB11 => MEM_RADDR_11_net, ADDRB10 => 
        MEM_RADDR_10_net, ADDRB9 => MEM_RADDR_9_net, ADDRB8 => 
        MEM_RADDR_8_net, ADDRB7 => MEM_RADDR_7_net, ADDRB6 => 
        MEM_RADDR_6_net, ADDRB5 => MEM_RADDR_5_net, ADDRB4 => 
        MEM_RADDR_4_net, ADDRB3 => MEM_RADDR_3_net, ADDRB2 => 
        MEM_RADDR_2_net, ADDRB1 => MEM_RADDR_1_net, ADDRB0 => 
        MEM_RADDR_0_net, DINA8 => ByteData_GND, DINA7 => 
        ByteData_GND, DINA6 => ByteData_GND, DINA5 => 
        ByteData_GND, DINA4 => ByteData_GND, DINA3 => 
        ByteData_GND, DINA2 => ByteData_GND, DINA1 => 
        ByteData_GND, DINA0 => data_reg_0, DINB8 => ByteData_GND, 
        DINB7 => ByteData_GND, DINB6 => ByteData_GND, DINB5 => 
        ByteData_GND, DINB4 => ByteData_GND, DINB3 => 
        ByteData_GND, DINB2 => ByteData_GND, DINB1 => 
        ByteData_GND, DINB0 => ByteData_GND, WIDTHA0 => 
        ByteData_GND, WIDTHA1 => ByteData_GND, WIDTHB0 => 
        ByteData_GND, WIDTHB1 => ByteData_GND, PIPEA => 
        ByteData_GND, PIPEB => ByteData_GND, WMODEA => 
        ByteData_GND, WMODEB => ByteData_GND, BLKA => MEMWENEG, 
        BLKB => MEMRENEG, WENA => ByteData_GND, WENB => 
        ByteData_VCC, CLKA => PLL_Test1_0_Sys_66M_Clk, CLKB => 
        PLL_Test1_0_Sys_66M_Clk, RESET => CMOS_DrvX_0_LVDSen, 
        DOUTA8 => RAM4K9_QXI_0_inst_DOUTA8, DOUTA7 => 
        RAM4K9_QXI_0_inst_DOUTA7, DOUTA6 => 
        RAM4K9_QXI_0_inst_DOUTA6, DOUTA5 => 
        RAM4K9_QXI_0_inst_DOUTA5, DOUTA4 => 
        RAM4K9_QXI_0_inst_DOUTA4, DOUTA3 => 
        RAM4K9_QXI_0_inst_DOUTA3, DOUTA2 => 
        RAM4K9_QXI_0_inst_DOUTA2, DOUTA1 => 
        RAM4K9_QXI_0_inst_DOUTA1, DOUTA0 => RAM4K9_QXI_0_DOUTA0, 
        DOUTB8 => RAM4K9_QXI_0_inst_DOUTB8, DOUTB7 => 
        RAM4K9_QXI_0_inst_DOUTB7, DOUTB6 => 
        RAM4K9_QXI_0_inst_DOUTB6, DOUTB5 => 
        RAM4K9_QXI_0_inst_DOUTB5, DOUTB4 => 
        RAM4K9_QXI_0_inst_DOUTB4, DOUTB3 => 
        RAM4K9_QXI_0_inst_DOUTB3, DOUTB2 => 
        RAM4K9_QXI_0_inst_DOUTB2, DOUTB1 => 
        RAM4K9_QXI_0_inst_DOUTB1, DOUTB0 => QXI_0_net);
    
    AO1_10 : AO1
      port map(A => XOR2_0_Y, B => AO1_9_Y, C => AND2_52_Y, Y => 
        AO1_10_Y);
    
    XOR2_41 : XOR2
      port map(A => MEM_WADDR_9_net, B => ByteData_GND, Y => 
        XOR2_41_Y);
    
    XNOR2_24 : XNOR2
      port map(A => RBINNXTSHIFT_4_net, B => MEM_WADDR_4_net, Y
         => XNOR2_24_Y);
    
    DFN1P0_EMPTY : DFN1P0
      port map(D => EMPTYINT, CLK => PLL_Test1_0_Sys_66M_Clk, PRE
         => CMOS_DrvX_0_LVDSen, Q => \DFN1P0_EMPTY\);
    
    AO1_30 : AO1
      port map(A => XOR2_3_Y, B => AND2_15_Y, C => AND2_46_Y, Y
         => AO1_30_Y);
    
    AND2_41 : AND2
      port map(A => XOR2_50_Y, B => XOR2_7_Y, Y => AND2_41_Y);
    
    XOR2_69 : XOR2
      port map(A => MEM_WADDR_3_net, B => ByteData_GND, Y => 
        XOR2_69_Y);
    
    AO1_16 : AO1
      port map(A => AND2_48_Y, B => AO1_18_Y, C => AO1_32_Y, Y
         => AO1_16_Y);
    
    AND2_17 : AND2
      port map(A => XNOR2_23_Y, B => XNOR2_4_Y, Y => AND2_17_Y);
    
    XOR2_6 : XOR2
      port map(A => MEM_RADDR_1_net, B => ByteData_GND, Y => 
        XOR2_6_Y);
    
    AO1_29 : AO1
      port map(A => XOR2_60_Y, B => AO1_12_Y, C => AND2_2_Y, Y
         => AO1_29_Y);
    
    AO1_13 : AO1
      port map(A => AND2_43_Y, B => AO1_5_Y, C => AO1_28_Y, Y => 
        AO1_13_Y);
    
    AND2_54 : AND2
      port map(A => XOR2_16_Y, B => XOR2_66_Y, Y => AND2_54_Y);
    
    DFN1C0_MEM_WADDR_3_inst : DFN1C0
      port map(D => WBINNXTSHIFT_3_net, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => CMOS_DrvX_0_LVDSen_3, Q
         => MEM_WADDR_3_net);
    
    XOR2_53 : XOR2
      port map(A => MEM_RADDR_6_net, B => ByteData_GND, Y => 
        XOR2_53_Y);
    
    AO1_36 : AO1
      port map(A => XOR2_50_Y, B => AO1_16_Y, C => AND2_26_Y, Y
         => AO1_36_Y);
    
    XNOR2_23 : XNOR2
      port map(A => RBINNXTSHIFT_10_net, B => MEM_WADDR_10_net, Y
         => XNOR2_23_Y);
    
    DFN1C0_MEM_WADDR_12_inst : DFN1C0
      port map(D => WBINNXTSHIFT_12_net, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => CMOS_DrvX_0_LVDSen_3, Q
         => MEM_WADDR_12_net);
    
    AO1_33 : AO1
      port map(A => AND2_31_Y, B => AO1_8_Y, C => AO1_37_Y, Y => 
        AO1_33_Y);
    
    XOR2_12 : XOR2
      port map(A => MEM_WADDR_12_net, B => ByteData_GND, Y => 
        XOR2_12_Y);
    
    XNOR2_7 : XNOR2
      port map(A => RBINNXTSHIFT_1_net, B => MEM_WADDR_1_net, Y
         => XNOR2_7_Y);
    
    XNOR2_12 : XNOR2
      port map(A => RBINNXTSHIFT_0_net, B => MEM_WADDR_0_net, Y
         => XNOR2_12_Y);
    
    AND2_48 : AND2
      port map(A => XOR2_14_Y, B => XOR2_65_Y, Y => AND2_48_Y);
    
    AND2_45 : AND2
      port map(A => MEM_WADDR_1_net, B => ByteData_GND, Y => 
        AND2_45_Y);
    
    AO1_19 : AO1
      port map(A => XOR2_62_Y, B => AO1_25_Y, C => AND2_49_Y, Y
         => AO1_19_Y);
    
    DFN1C0_MEM_WADDR_11_inst : DFN1C0
      port map(D => WBINNXTSHIFT_11_net, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => CMOS_DrvX_0_LVDSen_3, Q
         => MEM_WADDR_11_net);
    
    AND2_59 : AND2
      port map(A => XOR2_62_Y, B => XOR2_58_Y, Y => AND2_59_Y);
    
    DFN1C0_MEM_RADDR_2_inst : DFN1C0
      port map(D => RBINNXTSHIFT_2_net, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => CMOS_DrvX_0_LVDSen_3, Q
         => MEM_RADDR_2_net);
    
    AND2_4 : AND2
      port map(A => MEM_RADDR_4_net, B => ByteData_GND, Y => 
        AND2_4_Y);
    
    AND2_FULLINT : AND2
      port map(A => AND3_1_Y, B => XOR2_40_Y, Y => FULLINT);
    
    DFN1C0_MEM_RADDR_1_inst : DFN1C0
      port map(D => RBINNXTSHIFT_1_net, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => CMOS_DrvX_0_LVDSen_3, Q
         => MEM_RADDR_1_net);
    
    XOR2_WBINNXTSHIFT_6_inst : XOR2
      port map(A => XOR2_59_Y, B => AO1_9_Y, Y => 
        WBINNXTSHIFT_6_net);
    
    XOR2_50 : XOR2
      port map(A => MEM_RADDR_10_net, B => ByteData_GND, Y => 
        XOR2_50_Y);
    
    XNOR2_5 : XNOR2
      port map(A => MEM_RADDR_5_net, B => WBINNXTSHIFT_5_net, Y
         => XNOR2_5_Y);
    
    AO1_5 : AO1
      port map(A => AND2_25_Y, B => AO1_25_Y, C => AO1_23_Y, Y
         => AO1_5_Y);
    
    XNOR2_16 : XNOR2
      port map(A => RBINNXTSHIFT_8_net, B => MEM_WADDR_8_net, Y
         => XNOR2_16_Y);
    
    RAM4K9_QXI_3_inst : RAM4K9
      port map(ADDRA11 => MEM_WADDR_11_net, ADDRA10 => 
        MEM_WADDR_10_net, ADDRA9 => MEM_WADDR_9_net, ADDRA8 => 
        MEM_WADDR_8_net, ADDRA7 => MEM_WADDR_7_net, ADDRA6 => 
        MEM_WADDR_6_net, ADDRA5 => MEM_WADDR_5_net, ADDRA4 => 
        MEM_WADDR_4_net, ADDRA3 => MEM_WADDR_3_net, ADDRA2 => 
        MEM_WADDR_2_net, ADDRA1 => MEM_WADDR_1_net, ADDRA0 => 
        MEM_WADDR_0_net, ADDRB11 => MEM_RADDR_11_net, ADDRB10 => 
        MEM_RADDR_10_net, ADDRB9 => MEM_RADDR_9_net, ADDRB8 => 
        MEM_RADDR_8_net, ADDRB7 => MEM_RADDR_7_net, ADDRB6 => 
        MEM_RADDR_6_net, ADDRB5 => MEM_RADDR_5_net, ADDRB4 => 
        MEM_RADDR_4_net, ADDRB3 => MEM_RADDR_3_net, ADDRB2 => 
        MEM_RADDR_2_net, ADDRB1 => MEM_RADDR_1_net, ADDRB0 => 
        MEM_RADDR_0_net, DINA8 => ByteData_GND, DINA7 => 
        ByteData_GND, DINA6 => ByteData_GND, DINA5 => 
        ByteData_GND, DINA4 => ByteData_GND, DINA3 => 
        ByteData_GND, DINA2 => ByteData_GND, DINA1 => 
        ByteData_GND, DINA0 => data_reg_2, DINB8 => ByteData_GND, 
        DINB7 => ByteData_GND, DINB6 => ByteData_GND, DINB5 => 
        ByteData_GND, DINB4 => ByteData_GND, DINB3 => 
        ByteData_GND, DINB2 => ByteData_GND, DINB1 => 
        ByteData_GND, DINB0 => ByteData_GND, WIDTHA0 => 
        ByteData_GND, WIDTHA1 => ByteData_GND, WIDTHB0 => 
        ByteData_GND, WIDTHB1 => ByteData_GND, PIPEA => 
        ByteData_GND, PIPEB => ByteData_GND, WMODEA => 
        ByteData_GND, WMODEB => ByteData_GND, BLKA => MEMWENEG, 
        BLKB => MEMRENEG, WENA => ByteData_GND, WENB => 
        ByteData_VCC, CLKA => PLL_Test1_0_Sys_66M_Clk, CLKB => 
        PLL_Test1_0_Sys_66M_Clk, RESET => CMOS_DrvX_0_LVDSen, 
        DOUTA8 => RAM4K9_QXI_3_inst_DOUTA8, DOUTA7 => 
        RAM4K9_QXI_3_inst_DOUTA7, DOUTA6 => 
        RAM4K9_QXI_3_inst_DOUTA6, DOUTA5 => 
        RAM4K9_QXI_3_inst_DOUTA5, DOUTA4 => 
        RAM4K9_QXI_3_inst_DOUTA4, DOUTA3 => 
        RAM4K9_QXI_3_inst_DOUTA3, DOUTA2 => 
        RAM4K9_QXI_3_inst_DOUTA2, DOUTA1 => 
        RAM4K9_QXI_3_inst_DOUTA1, DOUTA0 => RAM4K9_QXI_3_DOUTA0, 
        DOUTB8 => RAM4K9_QXI_3_inst_DOUTB8, DOUTB7 => 
        RAM4K9_QXI_3_inst_DOUTB7, DOUTB6 => 
        RAM4K9_QXI_3_inst_DOUTB6, DOUTB5 => 
        RAM4K9_QXI_3_inst_DOUTB5, DOUTB4 => 
        RAM4K9_QXI_3_inst_DOUTB4, DOUTB3 => 
        RAM4K9_QXI_3_inst_DOUTB3, DOUTB2 => 
        RAM4K9_QXI_3_inst_DOUTB2, DOUTB1 => 
        RAM4K9_QXI_3_inst_DOUTB1, DOUTB0 => QXI_3_net);
    
    XOR2_WBINNXTSHIFT_5_inst : XOR2
      port map(A => XOR2_38_Y, B => AO1_19_Y, Y => 
        WBINNXTSHIFT_5_net);
    
    AND2_8 : AND2
      port map(A => XOR2_19_Y, B => XOR2_41_Y, Y => AND2_8_Y);
    
    XOR2_3 : XOR2
      port map(A => MEM_RADDR_3_net, B => ByteData_GND, Y => 
        XOR2_3_Y);
    
    XOR2_51 : XOR2
      port map(A => MEM_RADDR_3_net, B => ByteData_GND, Y => 
        XOR2_51_Y);
    
    DFN1C0_MEM_RADDR_8_inst : DFN1C0
      port map(D => RBINNXTSHIFT_8_net, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => CMOS_DrvX_0_LVDSen_3, Q
         => MEM_RADDR_8_net);
    
    AO1_27 : AO1
      port map(A => XOR2_19_Y, B => AO1_5_Y, C => AND2_58_Y, Y
         => AO1_27_Y);
    
    XOR2_66 : XOR2
      port map(A => MEM_WADDR_3_net, B => ByteData_GND, Y => 
        XOR2_66_Y);
    
    AND2_56 : AND2
      port map(A => AND2_48_Y, B => AND2_41_Y, Y => AND2_56_Y);
    
    XOR2_RBINNXTSHIFT_6_inst : XOR2
      port map(A => XOR2_68_Y, B => AO1_2_Y, Y => 
        RBINNXTSHIFT_6_net);
    
    XOR2_73 : XOR2
      port map(A => MEM_RADDR_8_net, B => ByteData_GND, Y => 
        XOR2_73_Y);
    
    AND2_53 : AND2
      port map(A => XOR2_9_Y, B => XOR2_3_Y, Y => AND2_53_Y);
    
    AND3_7 : AND3
      port map(A => XNOR2_12_Y, B => XNOR2_7_Y, C => XNOR2_13_Y, 
        Y => AND3_7_Y);
    
    XOR2_RBINNXTSHIFT_12_inst : XOR2
      port map(A => XOR2_74_Y, B => AO1_34_Y, Y => 
        RBINNXTSHIFT_12_net);
    
    XOR2_RBINNXTSHIFT_11_inst : XOR2
      port map(A => XOR2_76_Y, B => AO1_36_Y, Y => 
        RBINNXTSHIFT_11_net);
    
    XOR2_RBINNXTSHIFT_5_inst : XOR2
      port map(A => XOR2_20_Y, B => AO1_11_Y, Y => 
        RBINNXTSHIFT_5_net);
    
    AO1_17 : AO1
      port map(A => XOR2_41_Y, B => AND2_58_Y, C => AND2_50_Y, Y
         => AO1_17_Y);
    
    XNOR2_17 : XNOR2
      port map(A => MEM_RADDR_1_net, B => WBINNXTSHIFT_1_net, Y
         => XNOR2_17_Y);
    
    AND3_4 : AND3
      port map(A => XNOR2_15_Y, B => XNOR2_8_Y, C => XNOR2_2_Y, Y
         => AND3_4_Y);
    
    DFN1C0_MEM_WADDR_7_inst : DFN1C0
      port map(D => WBINNXTSHIFT_7_net, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => CMOS_DrvX_0_LVDSen_3, Q
         => MEM_WADDR_7_net);
    
    RAM4K9_QXI_6_inst : RAM4K9
      port map(ADDRA11 => MEM_WADDR_11_net, ADDRA10 => 
        MEM_WADDR_10_net, ADDRA9 => MEM_WADDR_9_net, ADDRA8 => 
        MEM_WADDR_8_net, ADDRA7 => MEM_WADDR_7_net, ADDRA6 => 
        MEM_WADDR_6_net, ADDRA5 => MEM_WADDR_5_net, ADDRA4 => 
        MEM_WADDR_4_net, ADDRA3 => MEM_WADDR_3_net, ADDRA2 => 
        MEM_WADDR_2_net, ADDRA1 => MEM_WADDR_1_net, ADDRA0 => 
        MEM_WADDR_0_net, ADDRB11 => MEM_RADDR_11_net, ADDRB10 => 
        MEM_RADDR_10_net, ADDRB9 => MEM_RADDR_9_net, ADDRB8 => 
        MEM_RADDR_8_net, ADDRB7 => MEM_RADDR_7_net, ADDRB6 => 
        MEM_RADDR_6_net, ADDRB5 => MEM_RADDR_5_net, ADDRB4 => 
        MEM_RADDR_4_net, ADDRB3 => MEM_RADDR_3_net, ADDRB2 => 
        MEM_RADDR_2_net, ADDRB1 => MEM_RADDR_1_net, ADDRB0 => 
        MEM_RADDR_0_net, DINA8 => ByteData_GND, DINA7 => 
        ByteData_GND, DINA6 => ByteData_GND, DINA5 => 
        ByteData_GND, DINA4 => ByteData_GND, DINA3 => 
        ByteData_GND, DINA2 => ByteData_GND, DINA1 => 
        ByteData_GND, DINA0 => data_reg_6, DINB8 => ByteData_GND, 
        DINB7 => ByteData_GND, DINB6 => ByteData_GND, DINB5 => 
        ByteData_GND, DINB4 => ByteData_GND, DINB3 => 
        ByteData_GND, DINB2 => ByteData_GND, DINB1 => 
        ByteData_GND, DINB0 => ByteData_GND, WIDTHA0 => 
        ByteData_GND, WIDTHA1 => ByteData_GND, WIDTHB0 => 
        ByteData_GND, WIDTHB1 => ByteData_GND, PIPEA => 
        ByteData_GND, PIPEB => ByteData_GND, WMODEA => 
        ByteData_GND, WMODEB => ByteData_GND, BLKA => MEMWENEG, 
        BLKB => MEMRENEG, WENA => ByteData_GND, WENB => 
        ByteData_VCC, CLKA => PLL_Test1_0_Sys_66M_Clk, CLKB => 
        PLL_Test1_0_Sys_66M_Clk, RESET => CMOS_DrvX_0_LVDSen, 
        DOUTA8 => RAM4K9_QXI_6_inst_DOUTA8, DOUTA7 => 
        RAM4K9_QXI_6_inst_DOUTA7, DOUTA6 => 
        RAM4K9_QXI_6_inst_DOUTA6, DOUTA5 => 
        RAM4K9_QXI_6_inst_DOUTA5, DOUTA4 => 
        RAM4K9_QXI_6_inst_DOUTA4, DOUTA3 => 
        RAM4K9_QXI_6_inst_DOUTA3, DOUTA2 => 
        RAM4K9_QXI_6_inst_DOUTA2, DOUTA1 => 
        RAM4K9_QXI_6_inst_DOUTA1, DOUTA0 => RAM4K9_QXI_6_DOUTA0, 
        DOUTB8 => RAM4K9_QXI_6_inst_DOUTB8, DOUTB7 => 
        RAM4K9_QXI_6_inst_DOUTB7, DOUTB6 => 
        RAM4K9_QXI_6_inst_DOUTB6, DOUTB5 => 
        RAM4K9_QXI_6_inst_DOUTB5, DOUTB4 => 
        RAM4K9_QXI_6_inst_DOUTB4, DOUTB3 => 
        RAM4K9_QXI_6_inst_DOUTB3, DOUTB2 => 
        RAM4K9_QXI_6_inst_DOUTB2, DOUTB1 => 
        RAM4K9_QXI_6_inst_DOUTB1, DOUTB0 => QXI_6_net);
    
    AO1_37 : AO1
      port map(A => XOR2_4_Y, B => AND2_1_Y, C => AND2_30_Y, Y
         => AO1_37_Y);
    
    RAM4K9_QXI_2_inst : RAM4K9
      port map(ADDRA11 => MEM_WADDR_11_net, ADDRA10 => 
        MEM_WADDR_10_net, ADDRA9 => MEM_WADDR_9_net, ADDRA8 => 
        MEM_WADDR_8_net, ADDRA7 => MEM_WADDR_7_net, ADDRA6 => 
        MEM_WADDR_6_net, ADDRA5 => MEM_WADDR_5_net, ADDRA4 => 
        MEM_WADDR_4_net, ADDRA3 => MEM_WADDR_3_net, ADDRA2 => 
        MEM_WADDR_2_net, ADDRA1 => MEM_WADDR_1_net, ADDRA0 => 
        MEM_WADDR_0_net, ADDRB11 => MEM_RADDR_11_net, ADDRB10 => 
        MEM_RADDR_10_net, ADDRB9 => MEM_RADDR_9_net, ADDRB8 => 
        MEM_RADDR_8_net, ADDRB7 => MEM_RADDR_7_net, ADDRB6 => 
        MEM_RADDR_6_net, ADDRB5 => MEM_RADDR_5_net, ADDRB4 => 
        MEM_RADDR_4_net, ADDRB3 => MEM_RADDR_3_net, ADDRB2 => 
        MEM_RADDR_2_net, ADDRB1 => MEM_RADDR_1_net, ADDRB0 => 
        MEM_RADDR_0_net, DINA8 => ByteData_GND, DINA7 => 
        ByteData_GND, DINA6 => ByteData_GND, DINA5 => 
        ByteData_GND, DINA4 => ByteData_GND, DINA3 => 
        ByteData_GND, DINA2 => ByteData_GND, DINA1 => 
        ByteData_GND, DINA0 => data_reg_2, DINB8 => ByteData_GND, 
        DINB7 => ByteData_GND, DINB6 => ByteData_GND, DINB5 => 
        ByteData_GND, DINB4 => ByteData_GND, DINB3 => 
        ByteData_GND, DINB2 => ByteData_GND, DINB1 => 
        ByteData_GND, DINB0 => ByteData_GND, WIDTHA0 => 
        ByteData_GND, WIDTHA1 => ByteData_GND, WIDTHB0 => 
        ByteData_GND, WIDTHB1 => ByteData_GND, PIPEA => 
        ByteData_GND, PIPEB => ByteData_GND, WMODEA => 
        ByteData_GND, WMODEB => ByteData_GND, BLKA => MEMWENEG, 
        BLKB => MEMRENEG, WENA => ByteData_GND, WENB => 
        ByteData_VCC, CLKA => PLL_Test1_0_Sys_66M_Clk, CLKB => 
        PLL_Test1_0_Sys_66M_Clk, RESET => CMOS_DrvX_0_LVDSen, 
        DOUTA8 => RAM4K9_QXI_2_inst_DOUTA8, DOUTA7 => 
        RAM4K9_QXI_2_inst_DOUTA7, DOUTA6 => 
        RAM4K9_QXI_2_inst_DOUTA6, DOUTA5 => 
        RAM4K9_QXI_2_inst_DOUTA5, DOUTA4 => 
        RAM4K9_QXI_2_inst_DOUTA4, DOUTA3 => 
        RAM4K9_QXI_2_inst_DOUTA3, DOUTA2 => 
        RAM4K9_QXI_2_inst_DOUTA2, DOUTA1 => 
        RAM4K9_QXI_2_inst_DOUTA1, DOUTA0 => RAM4K9_QXI_2_DOUTA0, 
        DOUTB8 => RAM4K9_QXI_2_inst_DOUTB8, DOUTB7 => 
        RAM4K9_QXI_2_inst_DOUTB7, DOUTB6 => 
        RAM4K9_QXI_2_inst_DOUTB6, DOUTB5 => 
        RAM4K9_QXI_2_inst_DOUTB5, DOUTB4 => 
        RAM4K9_QXI_2_inst_DOUTB4, DOUTB3 => 
        RAM4K9_QXI_2_inst_DOUTB3, DOUTB2 => 
        RAM4K9_QXI_2_inst_DOUTB2, DOUTB1 => 
        RAM4K9_QXI_2_inst_DOUTB1, DOUTB0 => QXI_2_net);
    
    DFN1E1C0_Q_6_inst : DFN1E1C0
      port map(D => QXI_6_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => CMOS_DrvX_0_LVDSen, E => DVLDI, Q => Fifo_dout(6));
    
    XOR2_0 : XOR2
      port map(A => MEM_WADDR_6_net, B => ByteData_GND, Y => 
        XOR2_0_Y);
    
    NAND2_1 : NAND2
      port map(A => \DFN1P0_EMPTY\, B => ByteData_VCC, Y => 
        NAND2_1_Y);
    
    DFN1C0_MEM_RADDR_4_inst : DFN1C0
      port map(D => RBINNXTSHIFT_4_net, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => CMOS_DrvX_0_LVDSen_3, Q
         => MEM_RADDR_4_net);
    
    AO1_4 : AO1
      port map(A => XOR2_47_Y, B => AND2_52_Y, C => AND2_13_Y, Y
         => AO1_4_Y);
    
    XOR2_68 : XOR2
      port map(A => MEM_RADDR_6_net, B => ByteData_GND, Y => 
        XOR2_68_Y);
    
    DFN1C0_MEM_RADDR_9_inst : DFN1C0
      port map(D => RBINNXTSHIFT_9_net, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => CMOS_DrvX_0_LVDSen_3, Q
         => MEM_RADDR_9_net);
    
    XOR2_WBINNXTSHIFT_12_inst : XOR2
      port map(A => XOR2_12_Y, B => AO1_13_Y, Y => 
        WBINNXTSHIFT_12_net);
    
    XOR2_WBINNXTSHIFT_11_inst : XOR2
      port map(A => XOR2_49_Y, B => AO1_29_Y, Y => 
        WBINNXTSHIFT_11_net);
    
    XNOR2_14 : XNOR2
      port map(A => RBINNXTSHIFT_3_net, B => MEM_WADDR_3_net, Y
         => XNOR2_14_Y);
    
    RAM4K9_QXI_7_inst : RAM4K9
      port map(ADDRA11 => MEM_WADDR_11_net, ADDRA10 => 
        MEM_WADDR_10_net, ADDRA9 => MEM_WADDR_9_net, ADDRA8 => 
        MEM_WADDR_8_net, ADDRA7 => MEM_WADDR_7_net, ADDRA6 => 
        MEM_WADDR_6_net, ADDRA5 => MEM_WADDR_5_net, ADDRA4 => 
        MEM_WADDR_4_net, ADDRA3 => MEM_WADDR_3_net, ADDRA2 => 
        MEM_WADDR_2_net, ADDRA1 => MEM_WADDR_1_net, ADDRA0 => 
        MEM_WADDR_0_net, ADDRB11 => MEM_RADDR_11_net, ADDRB10 => 
        MEM_RADDR_10_net, ADDRB9 => MEM_RADDR_9_net, ADDRB8 => 
        MEM_RADDR_8_net, ADDRB7 => MEM_RADDR_7_net, ADDRB6 => 
        MEM_RADDR_6_net, ADDRB5 => MEM_RADDR_5_net, ADDRB4 => 
        MEM_RADDR_4_net, ADDRB3 => MEM_RADDR_3_net, ADDRB2 => 
        MEM_RADDR_2_net, ADDRB1 => MEM_RADDR_1_net, ADDRB0 => 
        MEM_RADDR_0_net, DINA8 => ByteData_GND, DINA7 => 
        ByteData_GND, DINA6 => ByteData_GND, DINA5 => 
        ByteData_GND, DINA4 => ByteData_GND, DINA3 => 
        ByteData_GND, DINA2 => ByteData_GND, DINA1 => 
        ByteData_GND, DINA0 => ByteData_GND, DINB8 => 
        ByteData_GND, DINB7 => ByteData_GND, DINB6 => 
        ByteData_GND, DINB5 => ByteData_GND, DINB4 => 
        ByteData_GND, DINB3 => ByteData_GND, DINB2 => 
        ByteData_GND, DINB1 => ByteData_GND, DINB0 => 
        ByteData_GND, WIDTHA0 => ByteData_GND, WIDTHA1 => 
        ByteData_GND, WIDTHB0 => ByteData_GND, WIDTHB1 => 
        ByteData_GND, PIPEA => ByteData_GND, PIPEB => 
        ByteData_GND, WMODEA => ByteData_GND, WMODEB => 
        ByteData_GND, BLKA => MEMWENEG, BLKB => MEMRENEG, WENA
         => ByteData_GND, WENB => ByteData_VCC, CLKA => 
        PLL_Test1_0_Sys_66M_Clk, CLKB => PLL_Test1_0_Sys_66M_Clk, 
        RESET => CMOS_DrvX_0_LVDSen, DOUTA8 => 
        RAM4K9_QXI_7_inst_DOUTA8, DOUTA7 => 
        RAM4K9_QXI_7_inst_DOUTA7, DOUTA6 => 
        RAM4K9_QXI_7_inst_DOUTA6, DOUTA5 => 
        RAM4K9_QXI_7_inst_DOUTA5, DOUTA4 => 
        RAM4K9_QXI_7_inst_DOUTA4, DOUTA3 => 
        RAM4K9_QXI_7_inst_DOUTA3, DOUTA2 => 
        RAM4K9_QXI_7_inst_DOUTA2, DOUTA1 => 
        RAM4K9_QXI_7_inst_DOUTA1, DOUTA0 => RAM4K9_QXI_7_DOUTA0, 
        DOUTB8 => RAM4K9_QXI_7_inst_DOUTB8, DOUTB7 => 
        RAM4K9_QXI_7_inst_DOUTB7, DOUTB6 => 
        RAM4K9_QXI_7_inst_DOUTB6, DOUTB5 => 
        RAM4K9_QXI_7_inst_DOUTB5, DOUTB4 => 
        RAM4K9_QXI_7_inst_DOUTB4, DOUTB3 => 
        RAM4K9_QXI_7_inst_DOUTB3, DOUTB2 => 
        RAM4K9_QXI_7_inst_DOUTB2, DOUTB1 => 
        RAM4K9_QXI_7_inst_DOUTB1, DOUTB0 => QXI_7_net);
    
    AO1_21 : AO1
      port map(A => XOR2_53_Y, B => AO1_2_Y, C => AND2_1_Y, Y => 
        AO1_21_Y);
    
    XOR2_36 : XOR2
      port map(A => MEM_RADDR_1_net, B => ByteData_GND, Y => 
        XOR2_36_Y);
    
    XOR2_74 : XOR2
      port map(A => MEM_RADDR_12_net, B => ByteData_GND, Y => 
        XOR2_74_Y);
    
    XNOR2_8 : XNOR2
      port map(A => MEM_RADDR_7_net, B => WBINNXTSHIFT_7_net, Y
         => XNOR2_8_Y);
    
    AND2_25 : AND2
      port map(A => AND2_59_Y, B => AND2_44_Y, Y => AND2_25_Y);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3;
use proasic3.all;

entity enc_8b10b is

    port( TenbitDout              : out   std_logic_vector(9 downto 0);
          Din_Delay4_6            : in    std_logic;
          Din_Delay4_5            : in    std_logic;
          Din_Delay4_7            : in    std_logic;
          Din_Delay4_2            : in    std_logic;
          Din_Delay4_0            : in    std_logic;
          Din_Delay4_1            : in    std_logic;
          CRC_Reg_6               : in    std_logic;
          CRC_Reg_5               : in    std_logic;
          CRC_Reg_7               : in    std_logic;
          CRC_Reg_2               : in    std_logic;
          CRC_Reg_0               : in    std_logic;
          CRC_Reg_1               : in    std_logic;
          Bit_En                  : in    std_logic;
          PLL_Test1_0_SysRst_O    : in    std_logic;
          PLL_Test1_0_Sys_66M_Clk : in    std_logic;
          Kin_Delay4              : in    std_logic;
          CRC_ResultAva           : in    std_logic;
          N_423                   : in    std_logic;
          N_422                   : in    std_logic;
          N_425                   : in    std_logic;
          N_426                   : in    std_logic
        );

end enc_8b10b;

architecture DEF_ARCH of enc_8b10b is 

  component OA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XNOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XNOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN0E1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AX1E
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO13
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component NOR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AX1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XO1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component XA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OAI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN0C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AO1D
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AO1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1D
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal NIO_1, \un4_nio\, un2_nio, nio, un2_s_1, un2_s_0, 
        \L31\, \un3_nd1s6_0\, \L13\, compls6_0_1, compls6_a4_1, 
        \LPDL4_RNIBSL81\, compls6_0_0, compls6_a3_1, compls6_a2_0, 
        compls6_a3_2, ND1S6_0_3, \ND1S6_a2\, \ND1S6_a1\, 
        ND1S6_0_0, \ND1S6_0_2\, ND1S6_a4_1, \ND1S6_a4_0\, 
        \ND1S6_a3\, \ND1S6_a0_2\, \ND1S6_a0_1\, \K4\, \L22_0_0\, 
        L22_0_tz, \un2_l31[0]_net_1\, compls6_a0_0, \LPDL4\, 
        compls6_a1_0, N_424, compls6_a4_0_0, pdl6_0, PD0S6, 
        \un7_l13_a1\, \un7_l13_a0\, \un1_l04_a1\, \un1_l04_a0\, 
        ND1S6_a3_0, compls6, N_1_i, \L31_0\, un1_l31, \un12_l31\, 
        \L22\, \L22_1\, NCO, un6_pd1s6, \L04\, SINT, SINT_tz_tz, 
        \H4\, ND1S4, DO_1, NDO, un3_compls6, EO_1, \un1_L13[0]\, 
        CO_1, BO_1, NBO, \l13\, \un2_l40_m3\, IO_1, \un1_L22[0]\, 
        \COMPLS6\, un7_l13, un21_l13, un1_l04, \l13_m2_e\, 
        \l13tt_m1_e\, \un2_l40_m2_e\, \un2_l40tt_m1_e\, \S\, 
        \un1_l13[0]_net_1\, N_421, N_427, N_428, \G4\, \F4\, 
        ND0S4, PD0S4, un1_njo, \GO_RNO_0\, PD1S4, \un2_pdl4_i[0]\, 
        \LPDL6\, PDL4, COMPLS4, FO_1, GO_1, HO_1, JO_1, \L40\, 
        \un14_l13\, \un1_pd1s6\, \un3_pd1s6[0]_net_1\, S_2, PDL6, 
        AO_1, \un1_PD0S6[0]\, \XLRESET\, \LRESET\, \GND\, \VCC\, 
        GND_0, VCC_0 : std_logic;

begin 


    LPDL4_RNIEOBH2 : OA1A
      port map(A => compls6_a4_1, B => N_425, C => 
        \LPDL4_RNIBSL81\, Y => compls6_0_1);
    
    un2_l40_m3 : MX2C
      port map(A => \un2_l40tt_m1_e\, B => \un2_l40_m2_e\, S => 
        CRC_ResultAva, Y => \un2_l40_m3\);
    
    ND1S6_a0_1 : NOR2B
      port map(A => N_424, B => N_426, Y => \ND1S6_a0_1\);
    
    LPDL4_RNIBC7O : OR3A
      port map(A => N_425, B => \LPDL4\, C => N_422, Y => 
        compls6_a3_2);
    
    L22_0_0 : OA1A
      port map(A => L22_0_tz, B => N_425, C => \un2_l31[0]_net_1\, 
        Y => \L22_0_0\);
    
    l13tt_m1_e : OR2A
      port map(A => Din_Delay4_0, B => Din_Delay4_1, Y => 
        \l13tt_m1_e\);
    
    IO_RNO_2 : OR2B
      port map(A => N_426, B => \L40\, Y => un2_nio);
    
    un2_l40tt_m1_e : NOR2B
      port map(A => Din_Delay4_1, B => Din_Delay4_0, Y => 
        \un2_l40tt_m1_e\);
    
    L13_0_tz : OA1
      port map(A => un7_l13, B => \l13\, C => N_424, Y => 
        L22_0_tz);
    
    K4_RNIRO4F1 : AOI1
      port map(A => \ND1S6_a0_2\, B => \ND1S6_a0_1\, C => \K4\, Y
         => ND1S6_0_0);
    
    DO_RNO : XOR3
      port map(A => compls6, B => NDO, C => un3_compls6, Y => 
        DO_1);
    
    BO_RNO : XNOR3
      port map(A => compls6, B => NBO, C => un3_compls6, Y => 
        BO_1);
    
    LPDL4_RNIC40G : NOR2A
      port map(A => N_422, B => \LPDL4\, Y => compls6_a0_0);
    
    K4_RNIRN7AR : MX2
      port map(A => PD0S6, B => \un3_pd1s6[0]_net_1\, S => 
        \COMPLS6\, Y => \un1_PD0S6[0]\);
    
    LPDL4_RNINSULB : XNOR2
      port map(A => un3_compls6, B => compls6, Y => \COMPLS6\);
    
    LPDL4_RNIIF96B1 : AO1B
      port map(A => pdl6_0, B => \un3_pd1s6[0]_net_1\, C => 
        \un1_PD0S6[0]\, Y => PDL6);
    
    un7_l13_a0 : OR3A
      port map(A => Din_Delay4_1, B => Din_Delay4_0, C => 
        CRC_ResultAva, Y => \un7_l13_a0\);
    
    L13 : AO1
      port map(A => N_425, B => L22_0_tz, C => \un1_l13[0]_net_1\, 
        Y => \L13\);
    
    DO : DFN0E1C0
      port map(D => DO_1, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        \LRESET\, E => Bit_En, Q => TenbitDout(3));
    
    BO : DFN0E1C0
      port map(D => BO_1, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        \LRESET\, E => Bit_En, Q => TenbitDout(1));
    
    L22_1 : OR2B
      port map(A => N_425, B => \L31_0\, Y => \L22_1\);
    
    JO_RNO : AX1E
      port map(A => SINT, B => un1_njo, C => COMPLS4, Y => JO_1);
    
    H4_RNO : MX2
      port map(A => Din_Delay4_7, B => CRC_Reg_7, S => 
        CRC_ResultAva, Y => N_421);
    
    \FNS.un2_s_0\ : NOR2
      port map(A => N_426, B => N_425, Y => un2_s_0);
    
    S_RNI85BD : OR2
      port map(A => \S\, B => \K4\, Y => SINT_tz_tz);
    
    L04 : OR3C
      port map(A => un1_l04, B => N_424, C => N_425, Y => \L04\);
    
    K4_RNILF0I : AO13
      port map(A => \G4\, B => \F4\, C => \K4\, Y => PD1S4);
    
    l13_m2_e : OR2A
      port map(A => CRC_Reg_0, B => CRC_Reg_1, Y => \l13_m2_e\);
    
    AO_RNO : XOR2
      port map(A => N_422, B => \COMPLS6\, Y => AO_1);
    
    un1_l04_a0 : OR3
      port map(A => Din_Delay4_1, B => Din_Delay4_0, C => 
        CRC_ResultAva, Y => \un1_l04_a0\);
    
    XLRESET : DFN1
      port map(D => PLL_Test1_0_SysRst_O, CLK => 
        PLL_Test1_0_Sys_66M_Clk, Q => \XLRESET\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    un7_l13_0 : OR2B
      port map(A => \un7_l13_a1\, B => \un7_l13_a0\, Y => un7_l13);
    
    un21_l13_0 : OR2A
      port map(A => un1_l04, B => N_424, Y => un21_l13);
    
    LPDL4_RNI44TG1 : OR3C
      port map(A => \ND1S6_a4_0\, B => compls6_a0_0, C => un2_s_0, 
        Y => N_1_i);
    
    EO_RNO : XOR3
      port map(A => compls6, B => \un1_L13[0]\, C => un3_compls6, 
        Y => EO_1);
    
    un12_l31 : NOR3A
      port map(A => N_425, B => \un2_l40_m3\, C => N_424, Y => 
        \un12_l31\);
    
    EO_RNO_0 : MX2C
      port map(A => \L13\, B => \un14_l13\, S => N_426, Y => 
        \un1_L13[0]\);
    
    S_RNO : MX2A
      port map(A => \un4_nio\, B => un2_s_1, S => PDL6, Y => S_2);
    
    K4_RNI1OUG3 : NOR3C
      port map(A => \ND1S6_a2\, B => \ND1S6_a1\, C => ND1S6_0_0, 
        Y => ND1S6_0_3);
    
    G4_RNIBUVB : NOR2B
      port map(A => \G4\, B => \F4\, Y => ND1S4);
    
    ND1S6_a1_0 : NOR2B
      port map(A => N_423, B => N_422, Y => ND1S6_a3_0);
    
    AO : DFN0E1C0
      port map(D => AO_1, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        \LRESET\, E => Bit_En, Q => TenbitDout(0));
    
    LPDL4_RNIBSL81 : OR3A
      port map(A => N_425, B => compls6_a1_0, C => compls6_a3_1, 
        Y => \LPDL4_RNIBSL81\);
    
    HO_RNO : XOR2
      port map(A => \H4\, B => COMPLS4, Y => HO_1);
    
    un2_l40_m2_e : NOR2B
      port map(A => CRC_Reg_1, B => CRC_Reg_0, Y => 
        \un2_l40_m2_e\);
    
    un1_l31_0 : NOR2A
      port map(A => un7_l13, B => N_424, Y => un1_l31);
    
    LPDL4_RNI5C4P1 : AO1
      port map(A => compls6_a3_1, B => compls6_a2_0, C => 
        compls6_a3_2, Y => compls6_0_0);
    
    F4 : DFN0
      port map(D => N_427, CLK => PLL_Test1_0_Sys_66M_Clk, Q => 
        \F4\);
    
    compls6_a1_1 : OR2A
      port map(A => N_424, B => N_426, Y => compls6_a3_1);
    
    un3_nd1s6_0 : OR2A
      port map(A => N_426, B => \L13\, Y => \un3_nd1s6_0\);
    
    ND1S6_a4_0 : NOR2A
      port map(A => N_423, B => N_424, Y => \ND1S6_a4_0\);
    
    LPDL4_RNO_0 : AX1C
      port map(A => \LPDL6\, B => PD0S4, C => ND0S4, Y => 
        \un2_pdl4_i[0]\);
    
    LPDL4_RNIN8DR5 : OR3C
      port map(A => compls6_0_0, B => N_1_i, C => compls6_0_1, Y
         => compls6);
    
    ND1S6_a3 : OR3B
      port map(A => ND1S6_a3_0, B => N_426, C => N_425, Y => 
        \ND1S6_a3\);
    
    L31 : NOR3
      port map(A => \L31_0\, B => un1_l31, C => \un12_l31\, Y => 
        \L31\);
    
    JO_RNO_0 : XO1A
      port map(A => \F4\, B => \G4\, C => \H4\, Y => un1_njo);
    
    CO_RNO_1 : OR3C
      port map(A => un1_l04, B => N_424, C => N_426, Y => 
        un6_pd1s6);
    
    LPDL4_RNIE40G : OR2
      port map(A => \LPDL4\, B => N_423, Y => compls6_a1_0);
    
    l13_m3 : MX2C
      port map(A => \l13tt_m1_e\, B => \l13_m2_e\, S => 
        CRC_ResultAva, Y => \l13\);
    
    JO : DFN1E1C0
      port map(D => JO_1, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        \LRESET\, E => Bit_En, Q => TenbitDout(9));
    
    GND_i : GND
      port map(Y => \GND\);
    
    CO_RNO_0 : OR3C
      port map(A => un6_pd1s6, B => N_424, C => \L04\, Y => NCO);
    
    H4_RNII30I : OR2B
      port map(A => ND1S4, B => \H4\, Y => PD0S4);
    
    FO : DFN1E1C0
      port map(D => FO_1, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        \LRESET\, E => Bit_En, Q => TenbitDout(6));
    
    compls6_a2_0_0 : OR2
      port map(A => N_423, B => N_426, Y => compls6_a2_0);
    
    un7_l13_a1 : OR3B
      port map(A => CRC_Reg_1, B => CRC_ResultAva, C => CRC_Reg_0, 
        Y => \un7_l13_a1\);
    
    \un1_l13[0]\ : XA1
      port map(A => N_424, B => N_425, C => un1_l04, Y => 
        \un1_l13[0]_net_1\);
    
    CO : DFN0E1C0
      port map(D => CO_1, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        \LRESET\, E => Bit_En, Q => TenbitDout(2));
    
    GO_RNO_0 : NOR2
      port map(A => \H4\, B => \F4\, Y => \GO_RNO_0\);
    
    IO_RNO_3 : OR2B
      port map(A => Kin_Delay4, B => \L22\, Y => nio);
    
    LPDL6_RNILAP51 : MX2A
      port map(A => PD1S4, B => ND1S4, S => \LPDL6\, Y => COMPLS4);
    
    LPDL4_RNO : OAI1
      port map(A => COMPLS4, B => PD0S4, C => \un2_pdl4_i[0]\, Y
         => PDL4);
    
    LPDL4_RNI4KE01 : NOR3A
      port map(A => compls6_a4_0_0, B => \LPDL4\, C => N_422, Y
         => compls6_a4_1);
    
    IO_RNO : AX1E
      port map(A => \un1_L22[0]\, B => NIO_1, C => \COMPLS6\, Y
         => IO_1);
    
    LRESET : DFN0
      port map(D => \XLRESET\, CLK => PLL_Test1_0_Sys_66M_Clk, Q
         => \LRESET\);
    
    un1_l04_a1 : OR3A
      port map(A => CRC_ResultAva, B => CRC_Reg_1, C => CRC_Reg_0, 
        Y => \un1_l04_a1\);
    
    ND1S6_0_2 : AOI1B
      port map(A => ND1S6_a4_1, B => \ND1S6_a4_0\, C => 
        \ND1S6_a3\, Y => \ND1S6_0_2\);
    
    G4_RNO : MX2
      port map(A => Din_Delay4_6, B => CRC_Reg_6, S => 
        CRC_ResultAva, Y => N_428);
    
    F4_RNO : MX2
      port map(A => Din_Delay4_5, B => CRC_Reg_5, S => 
        CRC_ResultAva, Y => N_427);
    
    un14_l13 : OR3B
      port map(A => un1_l04, B => N_424, C => N_425, Y => 
        \un14_l13\);
    
    ND1S6_a2_1 : NOR2A
      port map(A => N_426, B => N_425, Y => ND1S6_a4_1);
    
    IO : DFN0E1C0
      port map(D => IO_1, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        \LRESET\, E => Bit_En, Q => TenbitDout(5));
    
    un1_l04_0 : OR2B
      port map(A => \un1_l04_a1\, B => \un1_l04_a0\, Y => un1_l04);
    
    LPDL4_RNI0KHQ5 : AO1B
      port map(A => ND1S6_0_3, B => \ND1S6_0_2\, C => \LPDL4\, Y
         => un3_compls6);
    
    H4_RNIQ8BV : OR3C
      port map(A => SINT_tz_tz, B => \H4\, C => ND1S4, Y => SINT);
    
    compls6_a4_0 : NOR2A
      port map(A => N_424, B => N_423, Y => compls6_a4_0_0);
    
    K4 : DFN0
      port map(D => Kin_Delay4, CLK => PLL_Test1_0_Sys_66M_Clk, Q
         => \K4\);
    
    IO_RNO_1 : NOR3C
      port map(A => \un4_nio\, B => un2_nio, C => nio, Y => NIO_1);
    
    H4 : DFN0
      port map(D => N_421, CLK => PLL_Test1_0_Sys_66M_Clk, Q => 
        \H4\);
    
    \un3_pd1s6[0]\ : MX2
      port map(A => \un1_pd1s6\, B => \un14_l13\, S => N_426, Y
         => \un3_pd1s6[0]_net_1\);
    
    L40 : NOR3
      port map(A => \un2_l40_m3\, B => N_424, C => N_425, Y => 
        \L40\);
    
    IO_RNO_0 : MX2A
      port map(A => \L22\, B => \L04\, S => N_426, Y => 
        \un1_L22[0]\);
    
    L31_0 : MX2B
      port map(A => \l13\, B => \un2_l40_m3\, S => N_424, Y => 
        \L31_0\);
    
    LPDL4 : DFN0C0
      port map(D => PDL4, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        \LRESET\, Q => \LPDL4\);
    
    G4 : DFN0
      port map(D => N_428, CLK => PLL_Test1_0_Sys_66M_Clk, Q => 
        \G4\);
    
    \un2_l31[0]\ : MX2B
      port map(A => un21_l13, B => un1_l31, S => N_425, Y => 
        \un2_l31[0]_net_1\);
    
    un1_l31_m2 : MX2C
      port map(A => Din_Delay4_2, B => CRC_Reg_2, S => 
        CRC_ResultAva, Y => N_424);
    
    LPDL4_RNIJK3H7 : NOR2B
      port map(A => \LPDL4\, B => PD0S6, Y => pdl6_0);
    
    un1_pd1s6 : OR2A
      port map(A => \L31\, B => \L22\, Y => \un1_pd1s6\);
    
    un4_nio : OR3C
      port map(A => N_425, B => N_426, C => \L13\, Y => \un4_nio\);
    
    ND1S6_a2 : OR3B
      port map(A => N_422, B => ND1S6_a4_1, C => N_424, Y => 
        \ND1S6_a2\);
    
    HO : DFN1E1C0
      port map(D => HO_1, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        \LRESET\, E => Bit_En, Q => TenbitDout(8));
    
    EO : DFN0E1C0
      port map(D => EO_1, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        \LRESET\, E => Bit_En, Q => TenbitDout(4));
    
    DO_RNO_0 : AO1D
      port map(A => N_424, B => \un2_l40_m3\, C => N_425, Y => 
        NDO);
    
    ND1S6_a1 : OR3B
      port map(A => N_425, B => ND1S6_a3_0, C => N_424, Y => 
        \ND1S6_a1\);
    
    ND1S6_a0_2 : NOR3A
      port map(A => N_425, B => N_422, C => N_423, Y => 
        \ND1S6_a0_2\);
    
    LPDL6 : DFN1C0
      port map(D => PDL6, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        \LRESET\, Q => \LPDL6\);
    
    S_RNO_0 : NOR2A
      port map(A => un2_s_0, B => \L31\, Y => un2_s_1);
    
    S : DFN1C0
      port map(D => S_2, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        \LRESET\, Q => \S\);
    
    CO_RNO : XNOR3
      port map(A => compls6, B => NCO, C => un3_compls6, Y => 
        CO_1);
    
    BO_RNO_0 : AO1C
      port map(A => \L40\, B => N_423, C => \L04\, Y => NBO);
    
    L22 : OR2B
      port map(A => \L22_0_0\, B => \L22_1\, Y => \L22\);
    
    K4_RNI0OA97 : OA1B
      port map(A => \L22\, B => \un3_nd1s6_0\, C => \K4\, Y => 
        PD0S6);
    
    GO_RNO : AX1D
      port map(A => \G4\, B => \GO_RNO_0\, C => COMPLS4, Y => 
        GO_1);
    
    FO_RNO : AX1C
      port map(A => \F4\, B => SINT, C => COMPLS4, Y => FO_1);
    
    GO : DFN1E1C0
      port map(D => GO_1, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        \LRESET\, E => Bit_En, Q => TenbitDout(7));
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    LPDL4_RNO_1 : OR2
      port map(A => \G4\, B => \F4\, Y => ND0S4);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3;
use proasic3.all;

entity FrameMk is

    port( FrameMk_GND             : in    std_logic;
          CMOS_DrvX_0_LVDSen_3    : in    std_logic;
          FrameMk_VCC             : in    std_logic;
          CMOS_DrvX_0_LVDSen      : in    std_logic;
          tok_c                   : out   std_logic;
          LVDS_O_c                : out   std_logic;
          Main_ctl4SD_0_ByteRdEn  : in    std_logic;
          CMOS_DrvX_0_LVDSen_2    : in    std_logic;
          CMOS_DrvX_0_LVDSen_1    : in    std_logic;
          CMOS_DrvX_0_LVDSen_0    : in    std_logic;
          FrameMk_0_LVDS_ok       : out   std_logic;
          FrameMk_0_LVDS_ok_i     : out   std_logic;
          PLL_Test1_0_SysRst_O    : in    std_logic;
          PLL_Test1_0_Sys_66M_Clk : in    std_logic
        );

end FrameMk;

architecture DEF_ARCH of FrameMk is 

  component OR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E0C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AO1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XNOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OAI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1E
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component INV
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1D
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component OA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component WaveGenSingleZ19
    port( RE                      : out   std_logic;
          PLL_Test1_0_SysRst_O    : in    std_logic := 'U';
          PLL_Test1_0_Sys_66M_Clk : in    std_logic := 'U';
          REen                    : in    std_logic := 'U'
        );
  end component;

  component AO1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component ByteData
    port( Fifo_dout               : out   std_logic_vector(7 downto 0);
          data_reg_6              : in    std_logic := 'U';
          data_reg_0              : in    std_logic := 'U';
          data_reg_5              : in    std_logic := 'U';
          data_reg_2              : in    std_logic := 'U';
          WE                      : in    std_logic := 'U';
          RE                      : in    std_logic := 'U';
          CMOS_DrvX_0_LVDSen      : in    std_logic := 'U';
          ByteData_VCC            : in    std_logic := 'U';
          CMOS_DrvX_0_LVDSen_3    : in    std_logic := 'U';
          ByteData_GND            : in    std_logic := 'U';
          CMOS_DrvX_0_LVDSen_2    : in    std_logic := 'U';
          PLL_Test1_0_Sys_66M_Clk : in    std_logic := 'U'
        );
  end component;

  component AXOI4
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component enc_8b10b
    port( TenbitDout              : out   std_logic_vector(9 downto 0);
          Din_Delay4_6            : in    std_logic := 'U';
          Din_Delay4_5            : in    std_logic := 'U';
          Din_Delay4_7            : in    std_logic := 'U';
          Din_Delay4_2            : in    std_logic := 'U';
          Din_Delay4_0            : in    std_logic := 'U';
          Din_Delay4_1            : in    std_logic := 'U';
          CRC_Reg_6               : in    std_logic := 'U';
          CRC_Reg_5               : in    std_logic := 'U';
          CRC_Reg_7               : in    std_logic := 'U';
          CRC_Reg_2               : in    std_logic := 'U';
          CRC_Reg_0               : in    std_logic := 'U';
          CRC_Reg_1               : in    std_logic := 'U';
          Bit_En                  : in    std_logic := 'U';
          PLL_Test1_0_SysRst_O    : in    std_logic := 'U';
          PLL_Test1_0_Sys_66M_Clk : in    std_logic := 'U';
          Kin_Delay4              : in    std_logic := 'U';
          CRC_ResultAva           : in    std_logic := 'U';
          N_423                   : in    std_logic := 'U';
          N_422                   : in    std_logic := 'U';
          N_425                   : in    std_logic := 'U';
          N_426                   : in    std_logic := 'U'
        );
  end component;

  component AXOI5
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NAND2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

    signal \ClkEn_2\, clken2, \ClkEn_1\, \ClkEn_0\, N_329_0, 
        \Prstate[0]_net_1\, N_690_0, \StepCnt[3]_net_1\, N_692_0, 
        \CRC_ResultAva\, N_291_0, N_7, \ClkDivCnt[1]_net_1\, 
        \ClkDivCnt[0]_net_1\, StepCnt_n1_0_i_0_0, N_341, N_569, 
        N_6, un1_StepCnt_3_i_0, N_8, StepCnt_n2_0_i_0_0, 
        \StepCnt[0]_net_1\, \StepCnt[1]_net_1\, N_570, 
        \StepCnt[2]_net_1\, N_450, N_358, DataClkCnt_e11_0_0_0, 
        N_350, DataClkCnt_e11_0_0_a5_1_1, N_1004, 
        \CRC_Reg_14_2_i_1[14]\, \CRC_Reg[6]_net_1\, 
        \CRC_Reg_14_2_i_0[14]\, \CRC_Reg[13]_net_1\, 
        \CRC_Reg_14_2_i_1[21]\, \CRC_Reg_14_2_i_0[21]\, 
        \CRC_Reg[20]_net_1\, \CRC_Reg_14_2_i_1[29]\, 
        \CRC_Reg[21]_net_1\, \CRC_Reg_14_2_i_0[29]\, 
        \CRC_Reg[28]_net_1\, \CRC_Reg_14_2_i_1[37]\, 
        \CRC_Reg[29]_net_1\, \CRC_Reg_14_2_i_0[37]\, 
        \CRC_Reg[36]_net_1\, \CRC_Reg_14_2_i_1[38]\, 
        \CRC_Reg[30]_net_1\, \CRC_Reg_14_2_i_0[38]\, 
        \CRC_Reg[37]_net_1\, \CRC_Reg_14_2_i_1[39]\, 
        \CRC_Reg[31]_net_1\, \CRC_Reg_14_2_i_0[39]\, 
        \CRC_Reg[38]_net_1\, \CRC_Reg_14_2_i_0[31]\, 
        \CRC_Reg[23]_net_1\, \CRC_Reg_14_2_i_0[30]\, 
        \CRC_Reg[22]_net_1\, \CRC_Reg_14_2_i_0[20]\, 
        \CRC_Reg[12]_net_1\, \CRC_Reg_14_2_i_0[19]\, 
        \CRC_Reg[11]_net_1\, \CRC_Reg_14_i_0_1[28]\, 
        \CRC_Reg_14_i_0_0[28]\, \CRC_Reg[27]_net_1\, 
        \CRC_Reg_14_2_i_0[13]\, \CRC_Reg[5]_net_1\, 
        \CRC_Reg_14_2_i_0[12]\, \CRC_Reg[4]_net_1\, 
        \CRC_Reg_14_2_i_0[8]\, \CRC_Reg[0]_net_1\, 
        \CRC_Reg_14_2_i_0[22]\, \CRC_Reg_14_2_i_0[23]\, 
        \CRC_Reg_14_i_0_1[36]\, \CRC_Reg_14_i_0_0[36]\, 
        \CRC_Reg[35]_net_1\, \CRC_Reg_14_i_0_1[35]\, 
        \CRC_Reg_14_i_0_0[35]\, \CRC_Reg[34]_net_1\, 
        \CRC_Reg_14_i_0_0[34]\, \CRC_Reg[26]_net_1\, 
        \CRC_Reg_14_i_0_1[33]\, N_692, \CRC_Reg[25]_net_1\, 
        \CRC_Reg_14_i_0_0[33]\, \CRC_Reg[32]_net_1\, 
        \CRC_Reg_14_i_0_1[32]\, \CRC_Reg[24]_net_1\, 
        \CRC_Reg_14_i_0_0[32]\, \CRC_Reg_14_i_0_0[27]\, 
        \CRC_Reg_14_i_0_0[26]\, \CRC_Reg_14_i_0_1[25]\, 
        \CRC_Reg[17]_net_1\, \CRC_Reg_14_i_0_0[25]\, 
        \CRC_Reg_14_i_0_0[18]\, \CRC_Reg[10]_net_1\, 
        \CRC_Reg_14_i_0_0[17]\, \CRC_Reg[16]_net_1\, 
        \CRC_Reg_14_i_0_0[11]\, \CRC_Reg_14_i_0_0[10]\, 
        \CRC_Reg[2]_net_1\, \CRC_Reg_14_i_0_0[9]\, 
        \CRC_Reg[1]_net_1\, \CRC_Reg_14_2_i_0[24]\, 
        \CRC_Reg_14_2_i_0[16]\, \CRC_Reg[8]_net_1\, 
        \CRC_Reg_14_2_i_0[15]\, \CRC_Reg[7]_net_1\, 
        \DataClkCnt[10]_net_1\, \DataClkCnt[11]_net_1\, N_706_i, 
        \CRC_Reg_14_i_0_0[7]\, N_605, \CRC_Reg_14_i_0_0[6]\, 
        \ByteDout[6]_net_1\, N_609, \CRC_Reg_14_i_0_0[5]\, 
        \ByteDout[5]_net_1\, N_612, \CRC_Reg_14_i_0_1[4]\, N_614, 
        N_615, N_353, \CRC_Reg_14_i_0_1[3]\, N_617, N_618, 
        \CRC_Reg_14_i_0_1[2]\, N_620, N_621, 
        \CRC_Reg_14_i_0_1[1]\, N_623, N_624, \ByteDout_8_i_3[4]\, 
        N_705, \rowcnt[4]_net_1\, \ByteDout_8_i_1[4]\, 
        \ByteDout_8_i_2[4]\, \FrameCnt[0]_net_1\, N_709, N_335, 
        \ByteDout_RNO_4[4]_net_1\, \ByteDout_RNO_5[4]_net_1\, 
        N_1055, \ByteDout_8_i_2[5]\, \FrameCnt[1]_net_1\, 
        \ByteDout_RNO_5[5]_net_1\, \ByteDout_8_i_1[5]\, 
        \ByteDout_RNO_3[5]_net_1\, \ByteDout_RNO_4[5]_net_1\, 
        \ByteDout_8_i_1[3]\, \ByteDout_8_i_a5_2_1[3]\, N_693, 
        \ByteDout_8_i_0[3]\, \Prstate[4]_net_1\, \Fifo_dout[3]\, 
        N_1049, \ByteDout_8_i_0_3[2]\, \rowcnt[2]_net_1\, 
        \ByteDout_RNO_7[2]_net_1\, \ByteDout_8_i_0_1[2]\, N_633, 
        \ByteDout_RNO_4[2]_net_1\, \ByteDout_RNO_5[2]_net_1\, 
        \ByteDout_8_i_3[7]\, \FrameCnt[3]_net_1\, 
        \ByteDout_8_i_2[7]\, \ByteDout_RNO_3[7]_net_1\, 
        \ByteDout_8_i_0[7]\, N_708, \ByteDout_8_i_a5_0_0[7]\, 
        N_698, \ByteDout_RNO_6[7]_net_1\, \ByteDout_8_i_4[6]\, 
        \ByteDout_8_i_1[6]\, \ByteDout_8_i_2[6]\, 
        \DelayCnt[3]_net_1\, \ByteDout_RNO_8[6]_net_1\, N_1067, 
        \ByteDout_RNO_6[6]_net_1\, N_1068, \ByteDout_8_1_4[0]\, 
        \ByteDout_8_1_2[0]\, \ByteDout_8_1_1[0]\, N_1033, 
        \ByteDout_8_1_a5_2_1[0]\, N_691, N_1037, N_1034, N_1035, 
        N_774, DataClkCnt_e2_i_0_0, N_298, \DataClkCnt[2]_net_1\, 
        DataClkCnt_e3_i_0_0, N_302, \DataClkCnt[3]_net_1\, 
        DataClkCnt_e4_i_0_0, N_305, \DataClkCnt[4]_net_1\, 
        DataClkCnt_e5_i_0_0, N_309, \DataClkCnt[5]_net_1\, 
        DataClkCnt_e6_i_0_0, N_314, \DataClkCnt[6]_net_1\, 
        \ByteDout_8_i_5[1]\, N_1047, \ByteDout_RNO_7[1]_net_1\, 
        N_1046, \ByteDout_8_i_2[1]\, \ByteDout_8_i_0[1]\, 
        \ByteDout_RNO_4[1]_net_1\, \ByteDout_RNO_5[1]_net_1\, 
        \Fifo_dout[1]\, N_1042, \Prstate_ns_i_0_0_a2_0[6]\, 
        \Prstate[1]_net_1\, DataClkCnt_e1_i_0_0, 
        \DataClkCnt[0]_net_1\, \DataClkCnt[1]_net_1\, 
        \ByteDout_8_i_0_a5_2_0[2]\, \DelayCnt[2]_net_1\, 
        \rowcnt[10]_net_1\, \PKGCnt[2]_net_1\, 
        DataClkCnt_e11_0_0_a5_0_0, \Prstate_ns_0_a5_0_2[3]\, 
        \Prstate_ns_0_a5_0_0[3]\, N_696, \Prstate[5]_net_1\, 
        \Prstate_ns_i_0_0_a5_0_0[2]\, \Prstate[6]_net_1\, 
        \Prstate_ns_0_a5_0_0[5]\, \Prstate[3]_net_1\, 
        \DelayCnt[1]_net_1\, \rowcnt[3]_net_1\, 
        \Prstate_ns_0_a5_1[0]\, N_368, CRC_ResultAva_3_0_a5_0, 
        \Prstate[7]_net_1\, \ByteDout_8_1_a5_3_0[0]\, 
        \PKGCnt[3]_net_1\, DelayCnt_c0, \Prstate_ns_0_a5_0[5]\, 
        \Prstate[2]_net_1\, \rowcnt[0]_net_1\, N_313, 
        CRC_ResultAva_3_0_o2_0, \ByteDout_8_i_0_a5_1_1[2]\, 
        DataOk_0_sqmuxa_0_a2_0_a5_9, \DataClkCnt[8]_net_1\, 
        DataOk_0_sqmuxa_0_a2_0_a5_6, \DataClkCnt[9]_net_1\, 
        DataOk_0_sqmuxa_0_a2_0_a5_8, \DataClkCnt[7]_net_1\, 
        DataOk_0_sqmuxa_0_a2_0_a5_4, DataOk_0_sqmuxa_0_a2_0_a5_7, 
        DataOk_0_sqmuxa_0_a2_0_a5_2, CRC_ResultAva_3_0_a5_0_2, 
        CRC_ResultAva_3_0_a5_0_1, clkdivcnt7_0, 
        \ClkDivCnt[3]_net_1\, \ClkDivCnt[2]_net_1\, clken2_0, 
        REen_1_0_0_a5_0, N_1126, N_333_i_0, DataClkCnt_e8, N_993, 
        N_994, N_995, N_290, N_443, N_688, N_288, N_442, N_686, 
        N_286, N_441, N_684, \CRC_Reg_RNO[9]_net_1\, N_440, N_682, 
        N_9, N_439, N_679, N_11, N_677, N_676, 
        \CRC_Reg_RNO[17]_net_1\, N_674, N_673, 
        \CRC_Reg_RNO[18]_net_1\, N_438, N_670, N_17, 
        \CRC_Reg_RNO[26]_net_1\, N_662, N_661, 
        \CRC_Reg_RNO[27]_net_1\, N_659, N_658, N_25, N_27, 
        \CRC_Reg[33]_net_1\, N_29, N_437, N_650, N_31, N_33, 
        N_261, N_642, N_641, N_259, N_639, N_638, N_12_i_0, 
        \ByteDout_RNO_1[2]_net_1\, N_256, N_436, N_629, N_254, 
        N_435, N_627, N_252, N_434, N_625, \CRC_Reg_RNO[1]_net_1\, 
        N_448, \CRC_Reg_RNO[2]_net_1\, \CRC_Reg_RNO[3]_net_1\, 
        \CRC_Reg[3]_net_1\, \CRC_Reg_RNO[4]_net_1\, 
        \CRC_Reg_RNO[5]_net_1\, N_610, \CRC_Reg_RNO[6]_net_1\, 
        N_607, \CRC_Reg_RNO[7]_net_1\, N_604, N_23, N_242, N_433, 
        N_599, N_240, N_432, N_597, N_238, N_431, N_595, N_236, 
        N_430, N_593, N_234, \CRC_Reg[39]_net_1\, N_232, N_230, 
        N_228, N_226, N_213, \CRC_Reg[14]_net_1\, N_186_i_0, 
        \ByteDout_RNO_1[7]_net_1\, N_184_i_0, 
        \ByteDout_RNO_0[6]_net_1\, \ByteDout_RNO_1[6]_net_1\, 
        N_182_i_0, \ByteDout_RNO_0[5]_net_1\, N_180_i_0, 
        \ByteDout_RNO_1[4]_net_1\, N_178_i_0, 
        \ByteDout_RNO_0[3]_net_1\, \ByteDout_RNO_2[3]_net_1\, 
        N_176_i_0, N_1045, \ByteDout_8[0]\, \PKGCnt[11]_net_1\, 
        N_1079_i, N_970, \CRC_Reg_RNO[0]_net_1\, N_577, N_576, 
        \Prstate_ns[0]\, \Prstate_RNO[1]_net_1\, N_1015, 
        DataClkCnt_e11, N_363, \PKGCnt[1]_net_1\, N_704, 
        \PKGCnt[0]_net_1\, \FrameCnt[8]_net_1\, N_381, 
        \PKGCnt[4]_net_1\, \PKGCnt[12]_net_1\, \rowcnt[9]_net_1\, 
        N_376, N_412, N_1030, N_5, N_323, \Prstate_RNO[3]_net_1\, 
        N_1084, N_548, DataOk_0_sqmuxa, N_997, N_330, N_999, 
        N_1001, DataClkCnt_e9, N_998, N_28, N_979, N_990, N_992, 
        N_26, N_24, N_22, N_20, N_18, N_16_i_0, N_1082, N_355, 
        N_150, N_1019, N_148, N_1017, \Prstate_RNO[5]_net_1\, 
        N_1012, N_1014, N_356, pts_en2, bit_en2, bit_en2_1, 
        data_reg27, \ByteSel[1]_net_1\, \ByteSel[2]_net_1\, 
        \ByteSel[0]_net_1\, data_reg28, \ByteDout_8_i_a5_4_0[1]\, 
        \ByteDout_8_i_a5_3_0[1]\, N_2220_tz, \FrameCnt[6]_net_1\, 
        \ByteDout_8_i_0_a5_0[2]\, ByteSel_n2, data_reg30, 
        ByteSel_1_sqmuxa, \Prstate_ns[7]\, 
        \Prstate_RNO_0[0]_net_1\, \PKGCnt[13]_net_1\, 
        \rowcnt[1]_net_1\, data_reg32, ByteSel_n0, ByteSel_n1, 
        N_721, N_414, N_702, \PKGCnt[6]_net_1\, \Fifo_dout[4]\, 
        \PKGCnt[15]_net_1\, \PKGCnt[7]_net_1\, \Fifo_dout[5]\, 
        \rowcnt[5]_net_1\, \PKGCnt[8]_net_1\, \Fifo_dout[6]\, 
        \PKGCnt[9]_net_1\, \rowcnt[6]_net_1\, \FrameCnt[2]_net_1\, 
        \Fifo_dout[7]\, \rowcnt[7]_net_1\, \ByteDout[0]_net_1\, 
        \CRC_Reg[19]_net_1\, \ByteDout[7]_net_1\, 
        \ByteDout[4]_net_1\, N_690, \ByteDout[3]_net_1\, 
        \ByteDout[2]_net_1\, \ByteDout[1]_net_1\, N_291, 
        \Fifo_dout[2]\, \PKGCnt[5]_net_1\, \CRC_Reg[15]_net_1\, 
        \CRC_Reg[18]_net_1\, \CRC_Reg[9]_net_1\, CRC_ResultAva_3, 
        \FrameCnt[5]_net_1\, \FrameCnt[4]_net_1\, 
        \rowcnt[8]_net_1\, N_413, \PKGCnt[14]_net_1\, 
        \FrameCnt[7]_net_1\, N_422, \Din_Delay4[0]_net_1\, N_425, 
        \Din_Delay4[3]_net_1\, \Prstate_ns[5]\, un1_Prstate_3_i, 
        N_746, N_419, \Prstate_RNO[6]_net_1\, \Fifo_dout[0]\, 
        N_329, \Shifter_4[8]\, \Shifter[9]_net_1\, 
        \TenbitDout[8]\, \PtS_En\, N_426, \Din_Delay4[4]_net_1\, 
        N_423, \Din_Delay4[1]_net_1\, \Shifter_4[7]\, 
        \Shifter[8]_net_1\, \TenbitDout[7]\, \Shifter_4[6]\, 
        \Shifter[7]_net_1\, \TenbitDout[6]\, \Shifter_4[5]\, 
        \Shifter[6]_net_1\, \TenbitDout[5]\, \Shifter_4[4]\, 
        \Shifter[5]_net_1\, \TenbitDout[4]\, \Shifter_4[3]\, 
        \Shifter[4]_net_1\, \TenbitDout[3]\, \Shifter_4[2]\, 
        \Shifter[3]_net_1\, \TenbitDout[2]\, \Shifter_4[1]\, 
        \Shifter[2]_net_1\, \TenbitDout[1]\, \Shifter_4[0]\, 
        \Shifter[1]_net_1\, \TenbitDout[0]\, StepCnt_n0, N_211, 
        N_394_i_i_0, StepCnte, \DataOk\, N_318, DataClkCnt_e10, 
        N_7_0, \PKGCnt[10]_net_1\, PKGCnt_n9, N_316, PKGCnt_n10, 
        PKGCnt_n11, N_325, PKGCnt_n12, PKGCnt_n13, N_347, 
        \Prstate_ns[3]\, PKGCnt_n14, PKGCnt_n15, N_403, rowcnt_n9, 
        N_334, rowcnt_n10, \FrameCnt_RNO[0]_net_1\, N_365, N_295, 
        N_300, N_304, N_306, N_310, N_312, N_320, N_322, N_327, 
        N_354, N_362, N_385_i, N_386_i, N_387_i, N_389_i_i_0, 
        N_390_i_i_0, \FrameCnt_RNO[2]_net_1\, N_392_i_i_0, 
        \PKGCnt_RNO[2]_net_1\, \FrameCnt_RNO[3]_net_1\, 
        \rowcnt_RNO[3]_net_1\, N_397_i_i_0, 
        \FrameCnt_RNO[4]_net_1\, \rowcnt_RNO[4]_net_1\, 
        \PKGCnt_RNO[4]_net_1\, \FrameCnt_RNO[5]_net_1\, 
        N_406_i_i_0, \PKGCnt_RNO[5]_net_1\, N_415_i_i_0, 
        \rowcnt_RNO[6]_net_1\, N_417_i_i_0, 
        \FrameCnt_RNO[7]_net_1\, N_444_i_i_0, 
        \PKGCnt_RNO[7]_net_1\, N_446_i_i_0, \rowcnt_RNO[8]_net_1\, 
        N_449_i_i_0, N_398_i, N_188, N_146, REen_1, \REen\, 
        FrameCnt_0_sqmuxa, \ClkDivCnt_3[1]\, I_5, 
        \ClkDivCnt_3[3]\, I_13, \WE\, \data_reg[2]_net_1\, 
        \data_reg[0]_net_1\, \Bit_En\, \ClkEn\, 
        \Shifter[0]_net_1\, \FrameMk_0_LVDS_ok\, \Kin_Delay1\, 
        \Kin\, \Kin_Delay4\, \Kin_Delay3\, \Kin_Delay2\, 
        \Din_Delay3[0]_net_1\, \Din_Delay2[0]_net_1\, 
        \Din_Delay3[1]_net_1\, \Din_Delay2[1]_net_1\, 
        \Din_Delay3[2]_net_1\, \Din_Delay2[2]_net_1\, 
        \Din_Delay3[3]_net_1\, \Din_Delay2[3]_net_1\, 
        \Din_Delay3[4]_net_1\, \Din_Delay2[4]_net_1\, 
        \Din_Delay3[5]_net_1\, \Din_Delay2[5]_net_1\, 
        \Din_Delay3[6]_net_1\, \Din_Delay2[6]_net_1\, 
        \Din_Delay3[7]_net_1\, \Din_Delay2[7]_net_1\, 
        \Din_Delay1[0]_net_1\, \Din_Delay1[1]_net_1\, 
        \Din_Delay1[2]_net_1\, \Din_Delay1[3]_net_1\, 
        \Din_Delay1[4]_net_1\, \Din_Delay1[5]_net_1\, 
        \Din_Delay1[6]_net_1\, \Din_Delay1[7]_net_1\, 
        \Din_Delay4[2]_net_1\, \Din_Delay4[5]_net_1\, 
        \Din_Delay4[6]_net_1\, \Din_Delay4[7]_net_1\, I_4, I_9, 
        \TenbitDout[9]\, \data_reg[5]_net_1\, \data_reg[6]_net_1\, 
        N_4, RE, \GND\, \VCC\, GND_0, VCC_0 : std_logic;

    for all : WaveGenSingleZ19
	Use entity work.WaveGenSingleZ19(DEF_ARCH);
    for all : ByteData
	Use entity work.ByteData(DEF_ARCH);
    for all : enc_8b10b
	Use entity work.enc_8b10b(DEF_ARCH);
begin 

    FrameMk_0_LVDS_ok <= \FrameMk_0_LVDS_ok\;

    \DataClkCnt_RNO_2[9]\ : OR3
      port map(A => N_706_i, B => \DataClkCnt[9]_net_1\, C => 
        N_330, Y => N_999);
    
    \CRC_Reg_RNO_0[7]\ : AO1A
      port map(A => \CRC_Reg[6]_net_1\, B => N_690_0, C => N_605, 
        Y => \CRC_Reg_14_i_0_0[7]\);
    
    \CRC_Reg_RNO_1[4]\ : NOR2
      port map(A => N_450, B => \ByteDout[4]_net_1\, Y => N_614);
    
    \rowcnt[3]\ : DFN1E0C0
      port map(D => \rowcnt_RNO[3]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => N_329, Q => \rowcnt[3]_net_1\);
    
    \Prstate_RNO[7]\ : OR3C
      port map(A => N_1079_i, B => CMOS_DrvX_0_LVDSen_1, C => 
        N_329_0, Y => \Prstate_ns[0]\);
    
    \CRC_Reg[21]\ : DFN1C0
      port map(D => N_226, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \CRC_Reg[21]_net_1\);
    
    \CRC_Reg_RNO_1[28]\ : AO1C
      port map(A => \CRC_Reg[27]_net_1\, B => N_690_0, C => 
        CMOS_DrvX_0_LVDSen_0, Y => \CRC_Reg_14_i_0_0[28]\);
    
    \rowcnt_RNO[8]\ : AX1
      port map(A => N_322, B => \rowcnt[7]_net_1\, C => 
        \rowcnt[8]_net_1\, Y => \rowcnt_RNO[8]_net_1\);
    
    \rowcnt_RNO[5]\ : XNOR2
      port map(A => \rowcnt[5]_net_1\, B => N_312, Y => 
        N_406_i_i_0);
    
    \Din_Delay1[0]\ : DFN1E1C0
      port map(D => \ByteDout[0]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => \ClkEn_1\, Q => \Din_Delay1[0]_net_1\);
    
    \Shifter_RNO[3]\ : MX2
      port map(A => \Shifter[4]_net_1\, B => \TenbitDout[3]\, S
         => \PtS_En\, Y => \Shifter_4[3]\);
    
    \PKGCnt_RNO[1]\ : XOR2
      port map(A => \PKGCnt[1]_net_1\, B => \PKGCnt[0]_net_1\, Y
         => N_386_i);
    
    \DataClkCnt_RNI17B6[5]\ : NOR2B
      port map(A => \DataClkCnt[5]_net_1\, B => 
        \DataClkCnt[6]_net_1\, Y => DataOk_0_sqmuxa_0_a2_0_a5_2);
    
    \DelayCnt_RNI9RS7_0[1]\ : NOR2A
      port map(A => DelayCnt_c0, B => \DelayCnt[1]_net_1\, Y => 
        N_381);
    
    \rowcnt[5]\ : DFN1E0C0
      port map(D => N_406_i_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => N_329, Q => 
        \rowcnt[5]_net_1\);
    
    \CRC_Reg[35]\ : DFN1C0
      port map(D => N_31, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \CRC_Reg[35]_net_1\);
    
    \CRC_Reg_RNO_1[34]\ : OAI1
      port map(A => \CRC_Reg[26]_net_1\, B => N_692_0, C => 
        CMOS_DrvX_0_LVDSen_0, Y => \CRC_Reg_14_i_0_0[34]\);
    
    \ByteDout_RNO_2[0]\ : NOR3C
      port map(A => N_1034, B => N_1035, C => N_774, Y => 
        \ByteDout_8_1_1[0]\);
    
    \DataClkCnt_RNO_0[6]\ : AX1E
      port map(A => N_314, B => \ClkEn_0\, C => 
        \DataClkCnt[6]_net_1\, Y => DataClkCnt_e6_i_0_0);
    
    \Din_Delay4_RNI1878[4]\ : MX2
      port map(A => \Din_Delay4[4]_net_1\, B => 
        \CRC_Reg[36]_net_1\, S => \CRC_ResultAva\, Y => N_426);
    
    Kin_Delay4 : DFN1E1P0
      port map(D => \Kin_Delay3\, CLK => PLL_Test1_0_Sys_66M_Clk, 
        PRE => PLL_Test1_0_SysRst_O, E => \ClkEn\, Q => 
        \Kin_Delay4\);
    
    \DelayCnt_RNIA8AH[1]\ : NOR2
      port map(A => N_698, B => N_696, Y => N_708);
    
    CRC_ResultAva_RNO_4 : OR2A
      port map(A => \CRC_ResultAva\, B => \Prstate[7]_net_1\, Y
         => CRC_ResultAva_3_0_a5_0);
    
    un1_clkdivcnt_I_4 : INV
      port map(A => \ClkDivCnt[0]_net_1\, Y => I_4);
    
    \StepCnt_RNO[0]\ : NOR3B
      port map(A => CMOS_DrvX_0_LVDSen_2, B => N_450, C => 
        \StepCnt[0]_net_1\, Y => StepCnt_n0);
    
    \Prstate_RNO[5]\ : NOR3A
      port map(A => CMOS_DrvX_0_LVDSen_1, B => N_1012, C => 
        N_1014, Y => \Prstate_RNO[5]_net_1\);
    
    \CRC_Reg_RNO[23]\ : NOR3
      port map(A => \CRC_Reg_14_2_i_0[23]\, B => N_642, C => 
        N_641, Y => N_261);
    
    CRC_ResultAva_RNIQ5FH : OR2A
      port map(A => N_692_0, B => N_690_0, Y => N_291_0);
    
    \ByteDout_RNO_4[3]\ : NOR3B
      port map(A => \DelayCnt[1]_net_1\, B => \DelayCnt[2]_net_1\, 
        C => \rowcnt[3]_net_1\, Y => \ByteDout_8_i_a5_2_1[3]\);
    
    \rowcnt[8]\ : DFN1E0C0
      port map(D => \rowcnt_RNO[8]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => N_329, Q => \rowcnt[8]_net_1\);
    
    DataOk_RNI116C : NOR2B
      port map(A => \DataOk\, B => \ClkEn_1\, Y => N_355);
    
    \ByteSel_RNO[0]\ : NOR2A
      port map(A => ByteSel_1_sqmuxa, B => \ByteSel[0]_net_1\, Y
         => ByteSel_n0);
    
    \CRC_Reg_RNO_1[33]\ : AO1C
      port map(A => \CRC_Reg[32]_net_1\, B => N_690_0, C => 
        CMOS_DrvX_0_LVDSen_0, Y => \CRC_Reg_14_i_0_0[33]\);
    
    \ByteDout_RNO_4[2]\ : OR2A
      port map(A => \Prstate[4]_net_1\, B => \Fifo_dout[2]\, Y
         => \ByteDout_RNO_4[2]_net_1\);
    
    \PKGCnt[11]\ : DFN1E0C0
      port map(D => PKGCnt_n11, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => N_329_0, Q => 
        \PKGCnt[11]_net_1\);
    
    \DelayCnt_RNI2DD9[3]\ : OR2A
      port map(A => \DelayCnt[3]_net_1\, B => N_691, Y => N_774);
    
    \CRC_Reg_RNO_1[30]\ : OAI1
      port map(A => \CRC_Reg[22]_net_1\, B => N_692_0, C => 
        CMOS_DrvX_0_LVDSen_0, Y => \CRC_Reg_14_2_i_0[30]\);
    
    ClkEn_1_RNI6E5E : OR2A
      port map(A => \ClkEn_1\, B => N_970, Y => N_450);
    
    \CRC_Reg_RNO_0[19]\ : XA1A
      port map(A => \CRC_Reg[39]_net_1\, B => \CRC_Reg[18]_net_1\, 
        C => N_690, Y => N_433);
    
    \CRC_Reg_RNO_1[18]\ : OAI1
      port map(A => \CRC_Reg[10]_net_1\, B => N_692, C => 
        CMOS_DrvX_0_LVDSen_1, Y => \CRC_Reg_14_i_0_0[18]\);
    
    \ClkDivCnt[1]\ : DFN1C0
      port map(D => \ClkDivCnt_3[1]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \ClkDivCnt[1]_net_1\);
    
    \CRC_Reg_RNO[29]\ : OA1B
      port map(A => \CRC_Reg[29]_net_1\, B => N_291_0, C => 
        \CRC_Reg_14_2_i_1[29]\, Y => N_228);
    
    \CRC_Reg[12]\ : DFN1C0
      port map(D => N_254, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \CRC_Reg[12]_net_1\);
    
    \Prstate_RNO_0[5]\ : AOI1
      port map(A => \Prstate[6]_net_1\, B => \ClkEn_0\, C => 
        \Prstate[5]_net_1\, Y => N_1012);
    
    \CRC_Reg_RNO_2[4]\ : NOR2A
      port map(A => N_690, B => \CRC_Reg[3]_net_1\, Y => N_615);
    
    \ByteSel[1]\ : DFN1C0
      port map(D => ByteSel_n1, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \ByteSel[1]_net_1\);
    
    \DelayCnt_RNIBRS7_0[1]\ : OR2
      port map(A => \DelayCnt[2]_net_1\, B => \DelayCnt[1]_net_1\, 
        Y => N_696);
    
    CRC_ResultAva_RNIHUQA : OR2B
      port map(A => \ClkEn_1\, B => \CRC_ResultAva\, Y => N_692);
    
    \Din_Delay2[7]\ : DFN1E1P0
      port map(D => \Din_Delay1[7]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, PRE => PLL_Test1_0_SysRst_O, E
         => \ClkEn_2\, Q => \Din_Delay2[7]_net_1\);
    
    \data_reg_RNO[2]\ : NOR2B
      port map(A => \ByteSel[2]_net_1\, B => \ByteSel[0]_net_1\, 
        Y => data_reg32);
    
    \CRC_Reg_RNO_0[24]\ : XA1A
      port map(A => \CRC_Reg[39]_net_1\, B => \CRC_Reg[23]_net_1\, 
        C => N_690, Y => N_441);
    
    \PKGCnt[6]\ : DFN1E0C0
      port map(D => N_417_i_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => N_329, Q => 
        \PKGCnt[6]_net_1\);
    
    \Prstate_RNIUUM8[7]\ : NOR2A
      port map(A => \ClkEn_0\, B => \Prstate[7]_net_1\, Y => 
        N_721);
    
    \PKGCnt_RNO_0[15]\ : OR3B
      port map(A => \PKGCnt[13]_net_1\, B => \PKGCnt[14]_net_1\, 
        C => N_347, Y => N_403);
    
    \Prstate_RNISS58[1]\ : NOR2
      port map(A => \Prstate[1]_net_1\, B => N_746, Y => 
        un1_Prstate_3_i);
    
    \CRC_Reg_RNO_2[19]\ : NOR2
      port map(A => N_291_0, B => \CRC_Reg[19]_net_1\, Y => N_599);
    
    \CRC_Reg[13]\ : DFN1C0
      port map(D => N_252, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \CRC_Reg[13]_net_1\);
    
    \CRC_Reg_RNO[14]\ : OA1B
      port map(A => \CRC_Reg[14]_net_1\, B => N_291_0, C => 
        \CRC_Reg_14_2_i_1[14]\, Y => N_213);
    
    \Prstate_RNO_0[0]\ : NOR2A
      port map(A => \Prstate[0]_net_1\, B => \ClkEn_0\, Y => 
        \Prstate_RNO_0[0]_net_1\);
    
    \DataClkCnt[2]\ : DFN1C0
      port map(D => N_18, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \DataClkCnt[2]_net_1\);
    
    \Prstate_RNO[3]\ : NOR3C
      port map(A => N_1084, B => CMOS_DrvX_0_LVDSen_1, C => N_548, 
        Y => \Prstate_RNO[3]_net_1\);
    
    \ClkDivCnt_RNIONNB[3]\ : OR2
      port map(A => \ClkDivCnt[3]_net_1\, B => 
        \ClkDivCnt[1]_net_1\, Y => clken2_0);
    
    \PKGCnt_RNO[13]\ : XNOR2
      port map(A => N_347, B => \PKGCnt[13]_net_1\, Y => 
        PKGCnt_n13);
    
    \Prstate_RNO[6]\ : NOR2A
      port map(A => CMOS_DrvX_0_LVDSen_2, B => N_419, Y => 
        \Prstate_RNO[6]_net_1\);
    
    \DataClkCnt_RNO_1[8]\ : OR2A
      port map(A => \DataClkCnt[8]_net_1\, B => \ClkEn_0\, Y => 
        N_994);
    
    \CRC_Reg_RNO_1[7]\ : NOR2
      port map(A => N_448, B => \CRC_Reg[7]_net_1\, Y => N_604);
    
    \CRC_Reg_RNO_0[23]\ : AO1C
      port map(A => \CRC_Reg[22]_net_1\, B => N_690_0, C => 
        CMOS_DrvX_0_LVDSen_0, Y => \CRC_Reg_14_2_i_0[23]\);
    
    \PKGCnt_RNO[7]\ : XOR2
      port map(A => \PKGCnt[7]_net_1\, B => N_306, Y => 
        \PKGCnt_RNO[7]_net_1\);
    
    \CRC_Reg_RNO_0[20]\ : XA1A
      port map(A => \CRC_Reg[39]_net_1\, B => \CRC_Reg[19]_net_1\, 
        C => N_690, Y => N_432);
    
    \Din_Delay4[3]\ : DFN1E1P0
      port map(D => \Din_Delay3[3]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, PRE => PLL_Test1_0_SysRst_O, E
         => \ClkEn\, Q => \Din_Delay4[3]_net_1\);
    
    \DataClkCnt_RNO_0[4]\ : AX1E
      port map(A => N_305, B => \ClkEn_0\, C => 
        \DataClkCnt[4]_net_1\, Y => DataClkCnt_e4_i_0_0);
    
    \CRC_Reg_RNO[5]\ : NOR3
      port map(A => N_353, B => \CRC_Reg_14_i_0_0[5]\, C => N_610, 
        Y => \CRC_Reg_RNO[5]_net_1\);
    
    \CRC_Reg[17]\ : DFN1C0
      port map(D => \CRC_Reg_RNO[17]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \CRC_Reg[17]_net_1\);
    
    \DataClkCnt_RNO[3]\ : NOR2A
      port map(A => N_979, B => DataClkCnt_e3_i_0_0, Y => N_20);
    
    \CRC_Reg_RNO[31]\ : NOR3
      port map(A => N_430, B => \CRC_Reg_14_2_i_0[31]\, C => 
        N_593, Y => N_236);
    
    \Prstate_RNIN2M8[0]\ : OR2B
      port map(A => \Prstate[0]_net_1\, B => \ClkEn_0\, Y => 
        N_329_0);
    
    PtS_En : DFN1C0
      port map(D => pts_en2, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \PtS_En\);
    
    \FrameCnt_RNO[1]\ : XOR2
      port map(A => \FrameCnt[1]_net_1\, B => \FrameCnt[0]_net_1\, 
        Y => N_387_i);
    
    \ByteDout_RNO_3[3]\ : NOR2A
      port map(A => N_413, B => \DelayCnt[2]_net_1\, Y => N_414);
    
    \PKGCnt[1]\ : DFN1E0C0
      port map(D => N_386_i, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => N_329_0, Q => 
        \PKGCnt[1]_net_1\);
    
    \Din_Delay1[5]\ : DFN1E1P0
      port map(D => \ByteDout[5]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, PRE => PLL_Test1_0_SysRst_O, E
         => \ClkEn_2\, Q => \Din_Delay1[5]_net_1\);
    
    \PKGCnt_RNO[12]\ : AX1C
      port map(A => N_325, B => \PKGCnt[11]_net_1\, C => 
        \PKGCnt[12]_net_1\, Y => PKGCnt_n12);
    
    \CRC_Reg[22]\ : DFN1C0
      port map(D => N_259, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \CRC_Reg[22]_net_1\);
    
    \CRC_Reg_RNO_1[8]\ : OAI1
      port map(A => \CRC_Reg[0]_net_1\, B => N_692_0, C => 
        CMOS_DrvX_0_LVDSen_0, Y => \CRC_Reg_14_2_i_0[8]\);
    
    \CRC_Reg_RNO[30]\ : NOR3
      port map(A => N_431, B => \CRC_Reg_14_2_i_0[30]\, C => 
        N_595, Y => N_238);
    
    \Shifter[6]\ : DFN1C0
      port map(D => \Shifter_4[6]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \Shifter[6]_net_1\);
    
    \DelayCnt_RNID8AH[1]\ : OR2
      port map(A => N_696, B => N_693, Y => N_702);
    
    \DataClkCnt_RNO_0[9]\ : OR3C
      port map(A => N_5, B => \DataClkCnt[9]_net_1\, C => N_330, 
        Y => N_997);
    
    \ByteDout_RNO_1[4]\ : OR3A
      port map(A => DelayCnt_c0, B => N_702, C => 
        \PKGCnt[7]_net_1\, Y => \ByteDout_RNO_1[4]_net_1\);
    
    \rowcnt_RNI39OD1[8]\ : OR3B
      port map(A => \rowcnt[7]_net_1\, B => \rowcnt[8]_net_1\, C
         => N_322, Y => N_334);
    
    \ByteSel_RNO[2]\ : XA1
      port map(A => \ByteSel[2]_net_1\, B => data_reg30, C => 
        ByteSel_1_sqmuxa, Y => ByteSel_n2);
    
    \rowcnt[10]\ : DFN1E0C0
      port map(D => rowcnt_n10, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => N_329, Q => 
        \rowcnt[10]_net_1\);
    
    \Din_Delay2[2]\ : DFN1E1P0
      port map(D => \Din_Delay1[2]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, PRE => PLL_Test1_0_SysRst_O, E
         => \ClkEn_2\, Q => \Din_Delay2[2]_net_1\);
    
    ClkEn_2 : DFN1C0
      port map(D => clken2, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \ClkEn_2\);
    
    \ByteDout_RNO_1[3]\ : OA1A
      port map(A => \ByteDout_8_i_a5_2_1[3]\, B => N_693, C => 
        \ByteDout_8_i_0[3]\, Y => \ByteDout_8_i_1[3]\);
    
    \ClkDivCnt_RNIE7FN[2]\ : NOR3
      port map(A => \ClkDivCnt[0]_net_1\, B => 
        \ClkDivCnt[2]_net_1\, C => clken2_0, Y => clken2);
    
    \Din_Delay1[7]\ : DFN1E1P0
      port map(D => \ByteDout[7]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, PRE => PLL_Test1_0_SysRst_O, E
         => \ClkEn_2\, Q => \Din_Delay1[7]_net_1\);
    
    PtS_En_RNO : NOR3A
      port map(A => \ClkDivCnt[1]_net_1\, B => 
        \ClkDivCnt[2]_net_1\, C => \ClkDivCnt[0]_net_1\, Y => 
        pts_en2);
    
    \CRC_Reg[23]\ : DFN1C0
      port map(D => N_261, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \CRC_Reg[23]_net_1\);
    
    \Din_Delay1[4]\ : DFN1E1P0
      port map(D => \ByteDout[4]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, PRE => PLL_Test1_0_SysRst_O, E
         => \ClkEn_2\, Q => \Din_Delay1[4]_net_1\);
    
    \Prstate_RNIV868_0[3]\ : NOR3
      port map(A => \Prstate[4]_net_1\, B => \Prstate[5]_net_1\, 
        C => \Prstate[3]_net_1\, Y => N_970);
    
    \CRC_Reg_RNO_0[2]\ : OR3
      port map(A => N_620, B => N_621, C => N_353, Y => 
        \CRC_Reg_14_i_0_1[2]\);
    
    \PKGCnt_RNI4DL91[7]\ : OR2B
      port map(A => \PKGCnt[7]_net_1\, B => N_306, Y => N_310);
    
    \CRC_Reg_RNO_0[9]\ : XA1A
      port map(A => \CRC_Reg[39]_net_1\, B => \CRC_Reg[8]_net_1\, 
        C => N_690, Y => N_440);
    
    \ByteDout_RNO_3[5]\ : OR3
      port map(A => N_704, B => \PKGCnt[0]_net_1\, C => N_698, Y
         => \ByteDout_RNO_3[5]_net_1\);
    
    \CRC_Reg_RNO_2[3]\ : NOR2A
      port map(A => N_690, B => \CRC_Reg[2]_net_1\, Y => N_618);
    
    \DataClkCnt_RNO_0[1]\ : AX1C
      port map(A => \DataClkCnt[0]_net_1\, B => \ClkEn_0\, C => 
        \DataClkCnt[1]_net_1\, Y => DataClkCnt_e1_i_0_0);
    
    \DataClkCnt[6]\ : DFN1C0
      port map(D => N_26, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \DataClkCnt[6]_net_1\);
    
    \FrameCnt_RNO[7]\ : XOR2
      port map(A => N_354, B => \FrameCnt[7]_net_1\, Y => 
        \FrameCnt_RNO[7]_net_1\);
    
    \CRC_Reg_RNO[28]\ : OA1B
      port map(A => \CRC_Reg[28]_net_1\, B => N_291_0, C => 
        \CRC_Reg_14_i_0_1[28]\, Y => N_23);
    
    \CRC_Reg_RNO[22]\ : NOR3
      port map(A => \CRC_Reg_14_2_i_0[22]\, B => N_639, C => 
        N_638, Y => N_259);
    
    \DataClkCnt[4]\ : DFN1C0
      port map(D => N_22, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \DataClkCnt[4]_net_1\);
    
    \CRC_Reg[38]\ : DFN1C0
      port map(D => N_232, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \CRC_Reg[38]_net_1\);
    
    \PKGCnt_RNO[6]\ : AX1C
      port map(A => N_300, B => \PKGCnt[5]_net_1\, C => 
        \PKGCnt[6]_net_1\, Y => N_417_i_i_0);
    
    \CRC_Reg[27]\ : DFN1C0
      port map(D => \CRC_Reg_RNO[27]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \CRC_Reg[27]_net_1\);
    
    \ByteDout_RNO_1[1]\ : NOR3C
      port map(A => \ByteDout_8_i_0[1]\, B => 
        \ByteDout_RNO_4[1]_net_1\, C => \ByteDout_RNO_5[1]_net_1\, 
        Y => \ByteDout_8_i_2[1]\);
    
    \ByteDout_RNO_7[6]\ : OR3
      port map(A => \DelayCnt[2]_net_1\, B => \PKGCnt[1]_net_1\, 
        C => N_698, Y => N_1068);
    
    \CRC_Reg_RNO[33]\ : OA1B
      port map(A => \CRC_Reg[33]_net_1\, B => N_291_0, C => 
        \CRC_Reg_14_i_0_1[33]\, Y => N_27);
    
    \ByteDout_RNO_1[5]\ : NOR3B
      port map(A => \ByteDout_RNO_3[5]_net_1\, B => 
        \ByteDout_RNO_4[5]_net_1\, C => N_335, Y => 
        \ByteDout_8_i_1[5]\);
    
    \CRC_Reg_RNO_0[35]\ : AO1D
      port map(A => N_692_0, B => \CRC_Reg[27]_net_1\, C => 
        \CRC_Reg_14_i_0_0[35]\, Y => \CRC_Reg_14_i_0_1[35]\);
    
    \Prstate_RNO_0[6]\ : MX2C
      port map(A => \Prstate[6]_net_1\, B => \Prstate[7]_net_1\, 
        S => \ClkEn_0\, Y => N_419);
    
    \CRC_Reg_RNO_0[37]\ : AO1D
      port map(A => N_692_0, B => \CRC_Reg[29]_net_1\, C => 
        \CRC_Reg_14_2_i_0[37]\, Y => \CRC_Reg_14_2_i_1[37]\);
    
    \CRC_Reg_RNO_1[38]\ : AO1C
      port map(A => \CRC_Reg[37]_net_1\, B => N_690_0, C => 
        CMOS_DrvX_0_LVDSen_0, Y => \CRC_Reg_14_2_i_0[38]\);
    
    \FrameCnt[5]\ : DFN1E0C0
      port map(D => \FrameCnt_RNO[5]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => N_365, Q => \FrameCnt[5]_net_1\);
    
    \DataClkCnt_RNIEK29[1]\ : NOR3C
      port map(A => \DataClkCnt[2]_net_1\, B => 
        \DataClkCnt[1]_net_1\, C => \Prstate[4]_net_1\, Y => 
        DataOk_0_sqmuxa_0_a2_0_a5_6);
    
    \CRC_Reg_RNO_0[36]\ : AO1D
      port map(A => N_692_0, B => \CRC_Reg[28]_net_1\, C => 
        \CRC_Reg_14_i_0_0[36]\, Y => \CRC_Reg_14_i_0_1[36]\);
    
    CRC_ResultAva_RNO_2 : AO1A
      port map(A => N_313, B => CRC_ResultAva_3_0_o2_0, C => 
        CRC_ResultAva_3_0_a5_0, Y => N_1030);
    
    \Prstate_RNO_1[7]\ : NOR3
      port map(A => \Prstate[1]_net_1\, B => \Prstate[0]_net_1\, 
        C => N_368, Y => \Prstate_ns_0_a5_1[0]\);
    
    \CRC_Reg_RNO[39]\ : OA1B
      port map(A => \CRC_Reg[39]_net_1\, B => N_291_0, C => 
        \CRC_Reg_14_2_i_1[39]\, Y => N_234);
    
    \DataClkCnt[0]\ : DFN1C0
      port map(D => N_7_0, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \DataClkCnt[0]_net_1\);
    
    \DelayCnt_RNI9RS7[1]\ : OR2B
      port map(A => \DelayCnt[1]_net_1\, B => DelayCnt_c0, Y => 
        N_313);
    
    \ClkDivCnt[2]\ : DFN1C0
      port map(D => I_9, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \ClkDivCnt[2]_net_1\);
    
    \Shifter_RNO[5]\ : MX2
      port map(A => \Shifter[6]_net_1\, B => \TenbitDout[5]\, S
         => \PtS_En\, Y => \Shifter_4[5]\);
    
    \data_reg_RNO[6]\ : NOR3A
      port map(A => \ByteSel[0]_net_1\, B => \ByteSel[1]_net_1\, 
        C => \ByteSel[2]_net_1\, Y => data_reg28);
    
    \CRC_Reg_RNO_1[3]\ : NOR2
      port map(A => N_450, B => \ByteDout[3]_net_1\, Y => N_617);
    
    Bit_En_RNO : NOR3A
      port map(A => \ClkDivCnt[2]_net_1\, B => 
        \ClkDivCnt[3]_net_1\, C => bit_en2_1, Y => bit_en2);
    
    \PKGCnt_RNIVB1Q[4]\ : NOR3B
      port map(A => \PKGCnt[3]_net_1\, B => \PKGCnt[4]_net_1\, C
         => N_295, Y => N_300);
    
    \Din_Delay4_RNIV778[3]\ : MX2C
      port map(A => \Din_Delay4[3]_net_1\, B => 
        \CRC_Reg[35]_net_1\, S => \CRC_ResultAva\, Y => N_425);
    
    \Shifter[8]\ : DFN1C0
      port map(D => \Shifter_4[8]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \Shifter[8]_net_1\);
    
    \Din_Delay4[6]\ : DFN1E1C0
      port map(D => \Din_Delay3[6]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => \ClkEn\, Q => \Din_Delay4[6]_net_1\);
    
    \PKGCnt[0]\ : DFN1C0
      port map(D => N_390_i_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \PKGCnt[0]_net_1\);
    
    \FrameCnt_RNO[4]\ : AX1C
      port map(A => \FrameCnt[3]_net_1\, B => N_320, C => 
        \FrameCnt[4]_net_1\, Y => \FrameCnt_RNO[4]_net_1\);
    
    \CRC_Reg[14]\ : DFN1C0
      port map(D => N_213, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \CRC_Reg[14]_net_1\);
    
    \FrameCnt_RNO[8]\ : AX1C
      port map(A => \FrameCnt[7]_net_1\, B => N_354, C => 
        \FrameCnt[8]_net_1\, Y => N_446_i_i_0);
    
    \DataClkCnt_RNO_1[11]\ : OR3A
      port map(A => \DataClkCnt[10]_net_1\, B => 
        \DataClkCnt[11]_net_1\, C => N_706_i, Y => 
        DataClkCnt_e11_0_0_a5_1_1);
    
    \rowcnt_RNIB3RM1[10]\ : OR3B
      port map(A => \rowcnt[9]_net_1\, B => \rowcnt[10]_net_1\, C
         => N_334, Y => N_362);
    
    \CRC_Reg_RNO_0[31]\ : XA1A
      port map(A => \CRC_Reg[39]_net_1\, B => \CRC_Reg[30]_net_1\, 
        C => N_690, Y => N_430);
    
    \CRC_Reg[19]\ : DFN1C0
      port map(D => N_242, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \CRC_Reg[19]_net_1\);
    
    \DataClkCnt_RNO_0[10]\ : OR3
      port map(A => N_706_i, B => \DataClkCnt[10]_net_1\, C => 
        N_350, Y => N_1001);
    
    \PKGCnt_RNO[15]\ : XNOR2
      port map(A => N_403, B => \PKGCnt[15]_net_1\, Y => 
        PKGCnt_n15);
    
    \Prstate_RNI9FL6[1]\ : OR2A
      port map(A => \Prstate[1]_net_1\, B => \DelayCnt[3]_net_1\, 
        Y => \Prstate_ns_i_0_0_a2_0[6]\);
    
    \DelayCnt_RNO_0[3]\ : AX1E
      port map(A => \DelayCnt[2]_net_1\, B => N_333_i_0, C => 
        \DelayCnt[3]_net_1\, Y => N_398_i);
    
    \CRC_Reg_RNO_0[4]\ : OR3
      port map(A => N_614, B => N_615, C => N_353, Y => 
        \CRC_Reg_14_i_0_1[4]\);
    
    \ByteSel_RNO[1]\ : XA1
      port map(A => \ByteSel[1]_net_1\, B => \ByteSel[0]_net_1\, 
        C => ByteSel_1_sqmuxa, Y => ByteSel_n1);
    
    \CRC_Reg_RNO_0[15]\ : XA1A
      port map(A => \CRC_Reg[39]_net_1\, B => \CRC_Reg[14]_net_1\, 
        C => N_690, Y => N_443);
    
    \Prstate_RNO_0[4]\ : NOR3B
      port map(A => CMOS_DrvX_0_LVDSen_1, B => 
        \Prstate_ns_0_a5_0_0[3]\, C => N_696, Y => 
        \Prstate_ns_0_a5_0_2[3]\);
    
    \Prstate_RNIARE5[2]\ : OR2
      port map(A => \Prstate[6]_net_1\, B => \Prstate[2]_net_1\, 
        Y => N_368);
    
    StepCnt_n2_0_i_0 : NOR2
      port map(A => un1_StepCnt_3_i_0, B => StepCnt_n2_0_i_0_0, Y
         => N_8);
    
    \Din_Delay1[3]\ : DFN1E1P0
      port map(D => \ByteDout[3]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, PRE => PLL_Test1_0_SysRst_O, E
         => \ClkEn_2\, Q => \Din_Delay1[3]_net_1\);
    
    \CRC_Reg_RNO_0[17]\ : AO1C
      port map(A => \CRC_Reg[16]_net_1\, B => N_690_0, C => 
        CMOS_DrvX_0_LVDSen_1, Y => \CRC_Reg_14_i_0_0[17]\);
    
    \Shifter[4]\ : DFN1C0
      port map(D => \Shifter_4[4]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \Shifter[4]_net_1\);
    
    \CRC_Reg_RNO_0[28]\ : AO1D
      port map(A => N_692_0, B => \CRC_Reg[20]_net_1\, C => 
        \CRC_Reg_14_i_0_0[28]\, Y => \CRC_Reg_14_i_0_1[28]\);
    
    \Prstate[6]\ : DFN1C0
      port map(D => \Prstate_RNO[6]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \Prstate[6]_net_1\);
    
    \CRC_Reg[4]\ : DFN1C0
      port map(D => \CRC_Reg_RNO[4]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \CRC_Reg[4]_net_1\);
    
    \CRC_Reg[2]\ : DFN1C0
      port map(D => \CRC_Reg_RNO[2]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \CRC_Reg[2]_net_1\);
    
    \CRC_Reg_RNO_0[16]\ : XA1A
      port map(A => \CRC_Reg[39]_net_1\, B => \CRC_Reg[15]_net_1\, 
        C => N_690, Y => N_442);
    
    \DelayCnt_RNO[2]\ : XA1B
      port map(A => \DelayCnt[2]_net_1\, B => N_333_i_0, C => 
        N_1019, Y => N_150);
    
    \ByteDout_RNO_4[7]\ : OA1A
      port map(A => \ByteDout_8_i_a5_0_0[7]\, B => N_698, C => 
        \ByteDout_RNO_6[7]_net_1\, Y => \ByteDout_8_i_0[7]\);
    
    \StepCnt_RNI6EU1[2]\ : NOR2B
      port map(A => \StepCnt[2]_net_1\, B => N_341, Y => N_358);
    
    \ByteSel_RNILSND[1]\ : AOI1B
      port map(A => \ByteSel[2]_net_1\, B => \ByteSel[1]_net_1\, 
        C => Main_ctl4SD_0_ByteRdEn, Y => ByteSel_1_sqmuxa);
    
    Kin_Delay2 : DFN1E1P0
      port map(D => \Kin_Delay1\, CLK => PLL_Test1_0_Sys_66M_Clk, 
        PRE => PLL_Test1_0_SysRst_O, E => \ClkEn\, Q => 
        \Kin_Delay2\);
    
    \CRC_Reg_RNO_2[9]\ : NOR2
      port map(A => N_291, B => \CRC_Reg[9]_net_1\, Y => N_682);
    
    \CRC_Reg_RNO_2[7]\ : NOR2
      port map(A => N_450, B => \ByteDout[7]_net_1\, Y => N_605);
    
    \Shifter[0]\ : DFN1C0
      port map(D => \Shifter_4[0]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \Shifter[0]_net_1\);
    
    StepCnt_n1_0_i_0 : NOR2
      port map(A => un1_StepCnt_3_i_0, B => StepCnt_n1_0_i_0_0, Y
         => N_6);
    
    \Prstate[7]\ : DFN1P0
      port map(D => \Prstate_ns[0]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, PRE => PLL_Test1_0_SysRst_O, Q
         => \Prstate[7]_net_1\);
    
    \DataClkCnt_RNO[5]\ : NOR2A
      port map(A => N_979, B => DataClkCnt_e5_i_0_0, Y => N_24);
    
    \Prstate[3]\ : DFN1C0
      port map(D => \Prstate_RNO[3]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \Prstate[3]_net_1\);
    
    \Din_Delay4_RNIP778[0]\ : MX2
      port map(A => \Din_Delay4[0]_net_1\, B => 
        \CRC_Reg[32]_net_1\, S => \CRC_ResultAva\, Y => N_422);
    
    \CRC_Reg_RNO_2[15]\ : NOR2
      port map(A => N_291, B => \CRC_Reg[15]_net_1\, Y => N_688);
    
    \DataClkCnt_RNIR2OV[9]\ : OR2A
      port map(A => \DataClkCnt[9]_net_1\, B => N_330, Y => N_350);
    
    \CRC_Reg_RNO_2[17]\ : NOR2
      port map(A => N_291, B => \CRC_Reg[17]_net_1\, Y => N_673);
    
    \CRC_Reg[31]\ : DFN1C0
      port map(D => N_236, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \CRC_Reg[31]_net_1\);
    
    \CRC_Reg_RNO_1[5]\ : NOR2
      port map(A => N_448, B => \CRC_Reg[5]_net_1\, Y => N_610);
    
    \PKGCnt[14]\ : DFN1E0C0
      port map(D => PKGCnt_n14, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => N_329_0, Q => 
        \PKGCnt[14]_net_1\);
    
    \CRC_Reg_RNO_0[32]\ : AO1D
      port map(A => N_692, B => \CRC_Reg[24]_net_1\, C => 
        \CRC_Reg_14_i_0_0[32]\, Y => \CRC_Reg_14_i_0_1[32]\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \DataClkCnt[10]\ : DFN1C0
      port map(D => DataClkCnt_e10, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \DataClkCnt[10]_net_1\);
    
    \DataClkCnt_RNO_0[11]\ : OA1
      port map(A => N_350, B => DataClkCnt_e11_0_0_a5_1_1, C => 
        N_1004, Y => DataClkCnt_e11_0_0_0);
    
    \CRC_Reg_RNO_2[16]\ : NOR2
      port map(A => N_291, B => \CRC_Reg[16]_net_1\, Y => N_686);
    
    \CRC_Reg_RNO_1[9]\ : OAI1
      port map(A => \CRC_Reg[1]_net_1\, B => N_692, C => 
        CMOS_DrvX_0_LVDSen_1, Y => \CRC_Reg_14_i_0_0[9]\);
    
    \ByteDout_RNO_7[1]\ : AO1
      port map(A => \ByteDout_8_i_a5_4_0[1]\, B => 
        \ByteDout_8_i_a5_3_0[1]\, C => N_691, Y => 
        \ByteDout_RNO_7[1]_net_1\);
    
    \FrameCnt[4]\ : DFN1E0C0
      port map(D => \FrameCnt_RNO[4]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => N_365, Q => \FrameCnt[4]_net_1\);
    
    \PKGCnt_RNO[9]\ : XOR2
      port map(A => N_316, B => \PKGCnt[9]_net_1\, Y => PKGCnt_n9);
    
    REGEN : WaveGenSingleZ19
      port map(RE => RE, PLL_Test1_0_SysRst_O => 
        PLL_Test1_0_SysRst_O, PLL_Test1_0_Sys_66M_Clk => 
        PLL_Test1_0_Sys_66M_Clk, REen => \REen\);
    
    \CRC_Reg_RNO_0[11]\ : AO1C
      port map(A => \CRC_Reg[10]_net_1\, B => N_690_0, C => 
        CMOS_DrvX_0_LVDSen_1, Y => \CRC_Reg_14_i_0_0[11]\);
    
    \rowcnt[9]\ : DFN1E0C0
      port map(D => rowcnt_n9, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => N_329, Q => 
        \rowcnt[9]_net_1\);
    
    \StepCnt_RNO[3]\ : AO1B
      port map(A => N_450, B => N_394_i_i_0, C => 
        CMOS_DrvX_0_LVDSen_2, Y => N_211);
    
    ClkEn_1_RNI325E : NOR2B
      port map(A => un1_Prstate_3_i, B => \ClkEn_1\, Y => N_1019);
    
    un1_clkdivcnt_I_8 : NOR2B
      port map(A => \ClkDivCnt[1]_net_1\, B => 
        \ClkDivCnt[0]_net_1\, Y => N_7);
    
    \CRC_Reg_RNO[6]\ : NOR3
      port map(A => N_353, B => \CRC_Reg_14_i_0_0[6]\, C => N_607, 
        Y => \CRC_Reg_RNO[6]_net_1\);
    
    \CRC_Reg_RNO[27]\ : NOR3
      port map(A => \CRC_Reg_14_i_0_0[27]\, B => N_659, C => 
        N_658, Y => \CRC_Reg_RNO[27]_net_1\);
    
    \Din_Delay2[3]\ : DFN1E1P0
      port map(D => \Din_Delay1[3]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, PRE => PLL_Test1_0_SysRst_O, E
         => \ClkEn_2\, Q => \Din_Delay2[3]_net_1\);
    
    \CRC_Reg[24]\ : DFN1C0
      port map(D => N_286, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \CRC_Reg[24]_net_1\);
    
    \CRC_Reg[29]\ : DFN1C0
      port map(D => N_228, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \CRC_Reg[29]_net_1\);
    
    LVDS_ok : DFN1E1C0
      port map(D => FrameCnt_0_sqmuxa, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => \ClkEn\, Q => \FrameMk_0_LVDS_ok\);
    
    \CRC_Reg_RNO[11]\ : NOR3
      port map(A => \CRC_Reg_14_i_0_0[11]\, B => N_677, C => 
        N_676, Y => N_11);
    
    \Prstate_RNO_2[5]\ : OR2A
      port map(A => \DelayCnt[3]_net_1\, B => \Prstate[6]_net_1\, 
        Y => \Prstate_ns_i_0_0_a5_0_0[2]\);
    
    \FrameCnt[1]\ : DFN1E0C0
      port map(D => N_387_i, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => N_365, Q => 
        \FrameCnt[1]_net_1\);
    
    \DataClkCnt[11]\ : DFN1C0
      port map(D => DataClkCnt_e11, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \DataClkCnt[11]_net_1\);
    
    \ByteDout_RNO_4[0]\ : NOR3B
      port map(A => \DelayCnt[2]_net_1\, B => \rowcnt[0]_net_1\, 
        C => N_313, Y => \ByteDout_8_1_a5_2_1[0]\);
    
    \CRC_Reg_RNO_2[27]\ : NOR2
      port map(A => N_291, B => \CRC_Reg[27]_net_1\, Y => N_658);
    
    \Prstate_RNO_0[3]\ : AO1
      port map(A => \Prstate[4]_net_1\, B => N_355, C => 
        \Prstate[3]_net_1\, Y => N_1084);
    
    \ByteDout_RNO_0[4]\ : OA1B
      port map(A => \FrameCnt[0]_net_1\, B => N_709, C => N_335, 
        Y => \ByteDout_8_i_2[4]\);
    
    \FrameCnt[3]\ : DFN1E0C0
      port map(D => \FrameCnt_RNO[3]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => N_365, Q => \FrameCnt[3]_net_1\);
    
    \CRC_Reg_RNO_2[26]\ : NOR2
      port map(A => N_291, B => \CRC_Reg[26]_net_1\, Y => N_661);
    
    \CRC_Reg_RNO[10]\ : NOR3
      port map(A => N_439, B => \CRC_Reg_14_i_0_0[10]\, C => 
        N_679, Y => N_9);
    
    \CRC_Reg_RNO[38]\ : OA1B
      port map(A => \CRC_Reg[38]_net_1\, B => N_291_0, C => 
        \CRC_Reg_14_2_i_1[38]\, Y => N_232);
    
    \CRC_Reg_RNO_2[11]\ : NOR2
      port map(A => N_291, B => \CRC_Reg[11]_net_1\, Y => N_676);
    
    \CRC_Reg_RNO[32]\ : OA1B
      port map(A => \CRC_Reg[32]_net_1\, B => N_291_0, C => 
        \CRC_Reg_14_i_0_1[32]\, Y => N_25);
    
    \rowcnt[0]\ : DFN1C0
      port map(D => N_389_i_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \rowcnt[0]_net_1\);
    
    CRC_ResultAva_RNIGUQA : OR2B
      port map(A => \ClkEn_0\, B => \CRC_ResultAva\, Y => N_692_0);
    
    \Prstate_RNIARE5[3]\ : OR2
      port map(A => \Prstate[5]_net_1\, B => \Prstate[3]_net_1\, 
        Y => N_746);
    
    CRC_ResultAva_RNO : AO1B
      port map(A => CRC_ResultAva_3_0_a5_0_2, B => 
        CRC_ResultAva_3_0_a5_0_1, C => N_1030, Y => 
        CRC_ResultAva_3);
    
    GenFIFO_Byte : ByteData
      port map(Fifo_dout(7) => \Fifo_dout[7]\, Fifo_dout(6) => 
        \Fifo_dout[6]\, Fifo_dout(5) => \Fifo_dout[5]\, 
        Fifo_dout(4) => \Fifo_dout[4]\, Fifo_dout(3) => 
        \Fifo_dout[3]\, Fifo_dout(2) => \Fifo_dout[2]\, 
        Fifo_dout(1) => \Fifo_dout[1]\, Fifo_dout(0) => 
        \Fifo_dout[0]\, data_reg_6 => \data_reg[6]_net_1\, 
        data_reg_0 => \data_reg[0]_net_1\, data_reg_5 => 
        \data_reg[5]_net_1\, data_reg_2 => \data_reg[2]_net_1\, 
        WE => \WE\, RE => RE, CMOS_DrvX_0_LVDSen => 
        CMOS_DrvX_0_LVDSen, ByteData_VCC => FrameMk_VCC, 
        CMOS_DrvX_0_LVDSen_3 => CMOS_DrvX_0_LVDSen_3, 
        ByteData_GND => FrameMk_GND, CMOS_DrvX_0_LVDSen_2 => 
        CMOS_DrvX_0_LVDSen_2, PLL_Test1_0_Sys_66M_Clk => 
        PLL_Test1_0_Sys_66M_Clk);
    
    \DataClkCnt_RNO_0[7]\ : AOI1
      port map(A => N_318, B => \ClkEn_1\, C => 
        \DataClkCnt[7]_net_1\, Y => N_990);
    
    \ByteDout_RNO_6[1]\ : OR3A
      port map(A => N_381, B => \PKGCnt[4]_net_1\, C => N_693, Y
         => N_1047);
    
    \ByteDout_RNO_8[2]\ : NOR3
      port map(A => \Prstate[6]_net_1\, B => \Prstate[0]_net_1\, 
        C => \Prstate[1]_net_1\, Y => \ByteDout_8_i_0_a5_1_1[2]\);
    
    \CRC_Reg_RNO_0[12]\ : XA1A
      port map(A => \CRC_Reg[39]_net_1\, B => \CRC_Reg[11]_net_1\, 
        C => N_690, Y => N_435);
    
    \rowcnt[6]\ : DFN1E0C0
      port map(D => \rowcnt_RNO[6]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => N_329, Q => \rowcnt[6]_net_1\);
    
    ClkEn_0 : DFN1C0
      port map(D => clken2, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \ClkEn_0\);
    
    \Prstate_RNIBVE5[5]\ : OR2A
      port map(A => \Prstate[5]_net_1\, B => \Prstate[4]_net_1\, 
        Y => N_691);
    
    \PKGCnt_RNO[10]\ : AX1C
      port map(A => N_316, B => \PKGCnt[9]_net_1\, C => 
        \PKGCnt[10]_net_1\, Y => PKGCnt_n10);
    
    ClkEn_1_RNI5HDH1_0 : OR2A
      port map(A => \ClkEn_1\, B => N_5, Y => N_979);
    
    ClkEn_1_RNI0K5H2 : AO1B
      port map(A => N_350, B => N_5, C => \ClkEn_1\, Y => N_363);
    
    \StepCnt[2]\ : DFN1E1C0
      port map(D => N_8, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => StepCnte, Q => 
        \StepCnt[2]_net_1\);
    
    \rowcnt_RNO[6]\ : AX1
      port map(A => N_312, B => \rowcnt[5]_net_1\, C => 
        \rowcnt[6]_net_1\, Y => \rowcnt_RNO[6]_net_1\);
    
    \rowcnt_RNIDFDP[4]\ : OR3C
      port map(A => N_304, B => \rowcnt[3]_net_1\, C => 
        \rowcnt[4]_net_1\, Y => N_312);
    
    \Din_Delay2[1]\ : DFN1E1C0
      port map(D => \Din_Delay1[1]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => \ClkEn_2\, Q => \Din_Delay2[1]_net_1\);
    
    \ByteDout[6]\ : DFN1E1C0
      port map(D => N_184_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => N_721, Q => 
        \ByteDout[6]_net_1\);
    
    \Shifter[5]\ : DFN1C0
      port map(D => \Shifter_4[5]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \Shifter[5]_net_1\);
    
    \PKGCnt[7]\ : DFN1E0C0
      port map(D => \PKGCnt_RNO[7]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => N_329, Q => \PKGCnt[7]_net_1\);
    
    \CRC_Reg_RNO_2[12]\ : NOR2
      port map(A => N_291, B => \CRC_Reg[12]_net_1\, Y => N_627);
    
    \ByteDout_RNO_6[6]\ : OR2A
      port map(A => \Prstate[4]_net_1\, B => \Fifo_dout[6]\, Y
         => \ByteDout_RNO_6[6]_net_1\);
    
    \Prstate_RNIV868[3]\ : OR3A
      port map(A => \Prstate[3]_net_1\, B => \Prstate[4]_net_1\, 
        C => \Prstate[5]_net_1\, Y => N_1049);
    
    \ByteDout_RNO_2[2]\ : OA1
      port map(A => N_705, B => \rowcnt[2]_net_1\, C => 
        \ByteDout_RNO_7[2]_net_1\, Y => \ByteDout_8_i_0_3[2]\);
    
    \ByteDout_RNO_4[1]\ : OR3
      port map(A => N_691, B => N_376, C => N_704, Y => 
        \ByteDout_RNO_4[1]_net_1\);
    
    \CRC_Reg[10]\ : DFN1C0
      port map(D => N_9, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \CRC_Reg[10]_net_1\);
    
    \FrameCnt[7]\ : DFN1E0C0
      port map(D => \FrameCnt_RNO[7]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => N_365, Q => \FrameCnt[7]_net_1\);
    
    \ClkDivCnt[0]\ : DFN1C0
      port map(D => I_4, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \ClkDivCnt[0]_net_1\);
    
    \CRC_Reg_RNO[13]\ : NOR3
      port map(A => N_434, B => \CRC_Reg_14_2_i_0[13]\, C => 
        N_625, Y => N_252);
    
    \DelayCnt_RNIETFO[2]\ : NOR3B
      port map(A => \DelayCnt[2]_net_1\, B => N_333_i_0, C => 
        \Prstate_ns_i_0_0_a2_0[6]\, Y => N_1126);
    
    \PKGCnt[12]\ : DFN1E0C0
      port map(D => PKGCnt_n12, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => N_329_0, Q => 
        \PKGCnt[12]_net_1\);
    
    \Shifter[7]\ : DFN1C0
      port map(D => \Shifter_4[7]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \Shifter[7]_net_1\);
    
    \DataClkCnt_RNI7FIS[8]\ : OR2A
      port map(A => \DataClkCnt[8]_net_1\, B => N_323, Y => N_330);
    
    \FrameCnt_RNO[6]\ : AX1C
      port map(A => \FrameCnt[5]_net_1\, B => N_327, C => 
        \FrameCnt[6]_net_1\, Y => N_415_i_i_0);
    
    \PKGCnt_RNO[4]\ : AX1
      port map(A => N_295, B => \PKGCnt[3]_net_1\, C => 
        \PKGCnt[4]_net_1\, Y => \PKGCnt_RNO[4]_net_1\);
    
    \Prstate_RNO_0[7]\ : OR3B
      port map(A => \Prstate_ns_0_a5_1[0]\, B => N_970, C => 
        \ClkEn_0\, Y => N_1079_i);
    
    \Prstate_RNIUBEB1[4]\ : NOR2A
      port map(A => \Prstate[4]_net_1\, B => DataOk_0_sqmuxa, Y
         => N_5);
    
    \DelayCnt[0]\ : DFN1C0
      port map(D => N_146, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => DelayCnt_c0);
    
    \DataClkCnt_RNI8C96[11]\ : NOR2A
      port map(A => \DataClkCnt[11]_net_1\, B => 
        \DataClkCnt[0]_net_1\, Y => DataOk_0_sqmuxa_0_a2_0_a5_4);
    
    \CRC_Reg_RNO[19]\ : NOR3
      port map(A => N_433, B => \CRC_Reg_14_2_i_0[19]\, C => 
        N_599, Y => N_242);
    
    \CRC_Reg_RNO_2[22]\ : NOR2
      port map(A => N_291, B => \CRC_Reg[22]_net_1\, Y => N_638);
    
    \CRC_Reg[32]\ : DFN1C0
      port map(D => N_25, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \CRC_Reg[32]_net_1\);
    
    \rowcnt_RNO[0]\ : XNOR2
      port map(A => \rowcnt[0]_net_1\, B => N_329_0, Y => 
        N_389_i_i_0);
    
    \ByteDout_RNO_5[1]\ : OR2
      port map(A => N_774, B => N_381, Y => 
        \ByteDout_RNO_5[1]_net_1\);
    
    \CRC_Reg_RNO_1[2]\ : NOR2
      port map(A => N_450, B => \ByteDout[2]_net_1\, Y => N_620);
    
    \DataClkCnt_RNIKRCP[7]\ : OR2B
      port map(A => N_318, B => \DataClkCnt[7]_net_1\, Y => N_323);
    
    \CRC_Reg_RNO_0[8]\ : XA1A
      port map(A => \CRC_Reg[39]_net_1\, B => \CRC_Reg[7]_net_1\, 
        C => N_690, Y => N_436);
    
    \DataClkCnt_RNO_0[8]\ : OR3C
      port map(A => N_5, B => \DataClkCnt[8]_net_1\, C => N_323, 
        Y => N_993);
    
    \data_reg[2]\ : DFN1C0
      port map(D => data_reg32, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \data_reg[2]_net_1\);
    
    \DelayCnt_RNIVCD9[0]\ : OR2
      port map(A => N_691, B => DelayCnt_c0, Y => N_698);
    
    \DelayCnt[1]\ : DFN1C0
      port map(D => N_148, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \DelayCnt[1]_net_1\);
    
    \CRC_Reg_RNO_0[34]\ : XA1A
      port map(A => \CRC_Reg[39]_net_1\, B => \CRC_Reg[33]_net_1\, 
        C => N_690, Y => N_437);
    
    \ByteSel[2]\ : DFN1C0
      port map(D => ByteSel_n2, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \ByteSel[2]_net_1\);
    
    ClkEn_1 : DFN1C0
      port map(D => clken2, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \ClkEn_1\);
    
    \rowcnt_RNO[10]\ : AX1
      port map(A => N_334, B => \rowcnt[9]_net_1\, C => 
        \rowcnt[10]_net_1\, Y => rowcnt_n10);
    
    \DataClkCnt_RNO_1[9]\ : OR2A
      port map(A => \DataClkCnt[9]_net_1\, B => \ClkEn_1\, Y => 
        N_998);
    
    \CRC_Reg[33]\ : DFN1C0
      port map(D => N_27, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \CRC_Reg[33]_net_1\);
    
    \DataClkCnt_RNO[8]\ : OR3C
      port map(A => N_993, B => N_994, C => N_995, Y => 
        DataClkCnt_e8);
    
    \CRC_Reg_RNO_0[0]\ : NOR2
      port map(A => N_450, B => \ByteDout[0]_net_1\, Y => N_577);
    
    \Shifter[2]\ : DFN1C0
      port map(D => \Shifter_4[2]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \Shifter[2]_net_1\);
    
    \CRC_Reg_RNO[7]\ : NOR3
      port map(A => N_353, B => \CRC_Reg_14_i_0_0[7]\, C => N_604, 
        Y => \CRC_Reg_RNO[7]_net_1\);
    
    \PKGCnt[5]\ : DFN1E0C0
      port map(D => \PKGCnt_RNO[5]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => N_329_0, Q => \PKGCnt[5]_net_1\);
    
    \CRC_Reg_RNO_0[3]\ : OR3
      port map(A => N_617, B => N_618, C => N_353, Y => 
        \CRC_Reg_14_i_0_1[3]\);
    
    \ByteDout_RNO_3[2]\ : OR3A
      port map(A => \ByteDout_8_i_0_a5_1_1[2]\, B => 
        \Prstate[4]_net_1\, C => \Prstate[5]_net_1\, Y => N_633);
    
    \StepCnt[0]\ : DFN1E1C0
      port map(D => StepCnt_n0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => StepCnte, Q => 
        \StepCnt[0]_net_1\);
    
    \DataClkCnt[7]\ : DFN1C0
      port map(D => N_28, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \DataClkCnt[7]_net_1\);
    
    \ByteDout_RNO[2]\ : NOR3C
      port map(A => \ByteDout_8_i_0_1[2]\, B => 
        \ByteDout_RNO_1[2]_net_1\, C => \ByteDout_8_i_0_3[2]\, Y
         => N_12_i_0);
    
    \CRC_Reg_RNO[37]\ : OA1B
      port map(A => \CRC_Reg[37]_net_1\, B => N_291_0, C => 
        \CRC_Reg_14_2_i_1[37]\, Y => N_230);
    
    \CRC_Reg[20]\ : DFN1C0
      port map(D => N_240, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \CRC_Reg[20]_net_1\);
    
    \Din_Delay4[4]\ : DFN1E1P0
      port map(D => \Din_Delay3[4]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, PRE => PLL_Test1_0_SysRst_O, E
         => \ClkEn\, Q => \Din_Delay4[4]_net_1\);
    
    \ByteDout_RNO[7]\ : NOR3C
      port map(A => \ByteDout_8_i_2[7]\, B => 
        \ByteDout_RNO_1[7]_net_1\, C => \ByteDout_8_i_3[7]\, Y
         => N_186_i_0);
    
    \PKGCnt_RNO[0]\ : XNOR2
      port map(A => \PKGCnt[0]_net_1\, B => N_329_0, Y => 
        N_390_i_i_0);
    
    \CRC_Reg_RNO[3]\ : OA1B
      port map(A => \CRC_Reg[3]_net_1\, B => N_448, C => 
        \CRC_Reg_14_i_0_1[3]\, Y => \CRC_Reg_RNO[3]_net_1\);
    
    \Prstate_RNO_0[1]\ : AOI1
      port map(A => \Prstate[2]_net_1\, B => \ClkEn_0\, C => 
        \Prstate[1]_net_1\, Y => N_1015);
    
    \CRC_Reg_RNO_0[33]\ : AO1D
      port map(A => N_692, B => \CRC_Reg[25]_net_1\, C => 
        \CRC_Reg_14_i_0_0[33]\, Y => \CRC_Reg_14_i_0_1[33]\);
    
    \ByteDout_RNO[0]\ : AO1B
      port map(A => \PKGCnt[11]_net_1\, B => N_708, C => 
        \ByteDout_8_1_4[0]\, Y => \ByteDout_8[0]\);
    
    \CRC_Reg[37]\ : DFN1C0
      port map(D => N_230, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \CRC_Reg[37]_net_1\);
    
    \ByteDout_RNO_1[6]\ : OR2
      port map(A => N_709, B => \FrameCnt[2]_net_1\, Y => 
        \ByteDout_RNO_1[6]_net_1\);
    
    \CRC_Reg_RNO_0[30]\ : XA1A
      port map(A => \CRC_Reg[39]_net_1\, B => \CRC_Reg[29]_net_1\, 
        C => N_690, Y => N_431);
    
    \Din_Delay2[6]\ : DFN1E1C0
      port map(D => \Din_Delay1[6]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => \ClkEn_2\, Q => \Din_Delay2[6]_net_1\);
    
    \ByteDout_RNO_0[5]\ : OR3A
      port map(A => DelayCnt_c0, B => N_702, C => 
        \PKGCnt[8]_net_1\, Y => \ByteDout_RNO_0[5]_net_1\);
    
    \Shifter_RNO[0]\ : MX2
      port map(A => \Shifter[1]_net_1\, B => \TenbitDout[0]\, S
         => \PtS_En\, Y => \Shifter_4[0]\);
    
    \PKGCnt[10]\ : DFN1E0C0
      port map(D => PKGCnt_n10, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => N_329_0, Q => 
        \PKGCnt[10]_net_1\);
    
    \ByteDout_RNO_9[1]\ : OR3
      port map(A => \Prstate[4]_net_1\, B => \Prstate[5]_net_1\, 
        C => \Prstate[2]_net_1\, Y => N_1042);
    
    \ByteDout_RNO_3[7]\ : OR2
      port map(A => \PKGCnt[10]_net_1\, B => N_702, Y => 
        \ByteDout_RNO_3[7]_net_1\);
    
    \rowcnt_RNIO28F[2]\ : NOR3C
      port map(A => \rowcnt[0]_net_1\, B => \rowcnt[1]_net_1\, C
         => \rowcnt[2]_net_1\, Y => N_304);
    
    \FrameCnt_RNO[2]\ : AX1C
      port map(A => \FrameCnt[0]_net_1\, B => \FrameCnt[1]_net_1\, 
        C => \FrameCnt[2]_net_1\, Y => \FrameCnt_RNO[2]_net_1\);
    
    \PKGCnt[4]\ : DFN1E0C0
      port map(D => \PKGCnt_RNO[4]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => N_329_0, Q => \PKGCnt[4]_net_1\);
    
    \Prstate_RNI15KA[3]\ : NOR3A
      port map(A => \Prstate[3]_net_1\, B => \DelayCnt[2]_net_1\, 
        C => \DelayCnt[3]_net_1\, Y => \Prstate_ns_0_a5_0_0[5]\);
    
    \ByteDout_RNO_2[7]\ : OA1B
      port map(A => \FrameCnt[3]_net_1\, B => N_709, C => N_335, 
        Y => \ByteDout_8_i_3[7]\);
    
    \CRC_Reg_RNO_1[29]\ : AO1C
      port map(A => \CRC_Reg[28]_net_1\, B => N_690_0, C => 
        CMOS_DrvX_0_LVDSen_0, Y => \CRC_Reg_14_2_i_0[29]\);
    
    \CRC_Reg_RNO[0]\ : NOR3
      port map(A => N_577, B => N_576, C => N_353, Y => 
        \CRC_Reg_RNO[0]_net_1\);
    
    \CRC_Reg_RNO_0[14]\ : AO1D
      port map(A => N_692_0, B => \CRC_Reg[6]_net_1\, C => 
        \CRC_Reg_14_2_i_0[14]\, Y => \CRC_Reg_14_2_i_1[14]\);
    
    ClkEn_1_RNI5HDH1 : OR2B
      port map(A => N_5, B => \ClkEn_1\, Y => N_706_i);
    
    LVDS_ok_RNO : NOR2A
      port map(A => \Prstate[0]_net_1\, B => N_362, Y => 
        FrameCnt_0_sqmuxa);
    
    \ByteDout_RNO_9[2]\ : OR2A
      port map(A => \DelayCnt[2]_net_1\, B => \rowcnt[10]_net_1\, 
        Y => \ByteDout_8_i_0_a5_2_0[2]\);
    
    \DataClkCnt_RNO_0[5]\ : AX1E
      port map(A => N_309, B => \ClkEn_0\, C => 
        \DataClkCnt[5]_net_1\, Y => DataClkCnt_e5_i_0_0);
    
    \Din_Delay4[0]\ : DFN1E1C0
      port map(D => \Din_Delay3[0]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => \ClkEn\, Q => \Din_Delay4[0]_net_1\);
    
    \data_reg_RNO[0]\ : NOR3
      port map(A => \ByteSel[1]_net_1\, B => \ByteSel[2]_net_1\, 
        C => \ByteSel[0]_net_1\, Y => data_reg27);
    
    \DataClkCnt_RNO[2]\ : NOR2A
      port map(A => N_979, B => DataClkCnt_e2_i_0_0, Y => N_18);
    
    \FrameCnt_RNIPUTE[6]\ : NOR3C
      port map(A => \FrameCnt[5]_net_1\, B => N_327, C => 
        \FrameCnt[6]_net_1\, Y => N_354);
    
    \Din_Delay3[5]\ : DFN1E1P0
      port map(D => \Din_Delay2[5]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, PRE => PLL_Test1_0_SysRst_O, E
         => \ClkEn_2\, Q => \Din_Delay3[5]_net_1\);
    
    \data_reg[5]\ : DFN1C0
      port map(D => data_reg30, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \data_reg[5]_net_1\);
    
    \DataClkCnt_RNO_0[3]\ : AX1E
      port map(A => N_302, B => \ClkEn_0\, C => 
        \DataClkCnt[3]_net_1\, Y => DataClkCnt_e3_i_0_0);
    
    \Prstate[2]\ : DFN1C0
      port map(D => \Prstate_ns[5]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \Prstate[2]_net_1\);
    
    \Prstate[5]\ : DFN1C0
      port map(D => \Prstate_RNO[5]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \Prstate[5]_net_1\);
    
    \CRC_Reg_RNO_0[13]\ : XA1A
      port map(A => \CRC_Reg[39]_net_1\, B => \CRC_Reg[12]_net_1\, 
        C => N_690, Y => N_434);
    
    \CRC_Reg_RNO[18]\ : NOR3
      port map(A => N_438, B => \CRC_Reg_14_i_0_0[18]\, C => 
        N_670, Y => \CRC_Reg_RNO[18]_net_1\);
    
    \CRC_Reg_RNO[12]\ : NOR3
      port map(A => N_435, B => \CRC_Reg_14_2_i_0[12]\, C => 
        N_627, Y => N_254);
    
    \CRC_Reg_RNO_0[10]\ : XA1A
      port map(A => \CRC_Reg[39]_net_1\, B => \CRC_Reg[9]_net_1\, 
        C => N_690, Y => N_439);
    
    \PKGCnt[13]\ : DFN1E0C0
      port map(D => PKGCnt_n13, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => N_329_0, Q => 
        \PKGCnt[13]_net_1\);
    
    \DataClkCnt_RNILRDF[8]\ : NOR3B
      port map(A => \DataClkCnt[8]_net_1\, B => 
        DataOk_0_sqmuxa_0_a2_0_a5_6, C => \DataClkCnt[9]_net_1\, 
        Y => DataOk_0_sqmuxa_0_a2_0_a5_9);
    
    \CRC_Reg_RNO[26]\ : NOR3
      port map(A => \CRC_Reg_14_i_0_0[26]\, B => N_662, C => 
        N_661, Y => \CRC_Reg_RNO[26]_net_1\);
    
    \ByteDout_RNO_1[0]\ : OA1A
      port map(A => \ByteDout_8_1_a5_2_1[0]\, B => N_691, C => 
        N_1037, Y => \ByteDout_8_1_2[0]\);
    
    StepCnt_n1_0_i_0_a5 : NOR2
      port map(A => \StepCnt[0]_net_1\, B => \StepCnt[1]_net_1\, 
        Y => N_569);
    
    \DataClkCnt[5]\ : DFN1C0
      port map(D => N_24, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \DataClkCnt[5]_net_1\);
    
    \CRC_Reg_RNO_1[19]\ : OAI1
      port map(A => \CRC_Reg[11]_net_1\, B => N_692_0, C => 
        CMOS_DrvX_0_LVDSen_0, Y => \CRC_Reg_14_2_i_0[19]\);
    
    \ByteDout_RNO_8[1]\ : OR3
      port map(A => \DelayCnt[1]_net_1\, B => \PKGCnt[12]_net_1\, 
        C => N_698, Y => N_1046);
    
    \ByteDout_RNO_8[6]\ : OR2
      port map(A => \PKGCnt[9]_net_1\, B => N_702, Y => 
        \ByteDout_RNO_8[6]_net_1\);
    
    REen : DFN1E1C0
      port map(D => REen_1, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => \ClkEn\, Q => \REen\);
    
    \Din_Delay2[0]\ : DFN1E1C0
      port map(D => \Din_Delay1[0]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => \ClkEn_2\, Q => \Din_Delay2[0]_net_1\);
    
    \DataClkCnt_RNIUDMC[3]\ : NOR3C
      port map(A => \DataClkCnt[4]_net_1\, B => 
        \DataClkCnt[3]_net_1\, C => DataOk_0_sqmuxa_0_a2_0_a5_2, 
        Y => DataOk_0_sqmuxa_0_a2_0_a5_7);
    
    StepCnt_n1_0_i_0_RNO : OR2
      port map(A => N_341, B => N_569, Y => StepCnt_n1_0_i_0_0);
    
    \CRC_Reg_RNO_2[24]\ : NOR2
      port map(A => N_291, B => \CRC_Reg[24]_net_1\, Y => N_684);
    
    \CRC_Reg_RNO_2[13]\ : NOR2
      port map(A => N_291, B => \CRC_Reg[13]_net_1\, Y => N_625);
    
    \CRC_Reg_RNO_2[10]\ : NOR2
      port map(A => N_291, B => \CRC_Reg[10]_net_1\, Y => N_679);
    
    \CRC_Reg[5]\ : DFN1C0
      port map(D => \CRC_Reg_RNO[5]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \CRC_Reg[5]_net_1\);
    
    \ByteDout_RNO_12[1]\ : OR2A
      port map(A => \DelayCnt[2]_net_1\, B => \DelayCnt[1]_net_1\, 
        Y => \ByteDout_8_i_a5_3_0[1]\);
    
    \DelayCnt[2]\ : DFN1C0
      port map(D => N_150, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \DelayCnt[2]_net_1\);
    
    \ByteDout_RNO_0[1]\ : OR3A
      port map(A => \DelayCnt[2]_net_1\, B => \rowcnt[9]_net_1\, 
        C => N_698, Y => N_1045);
    
    \ByteDout_RNO_7[2]\ : OR3A
      port map(A => DelayCnt_c0, B => N_702, C => 
        \PKGCnt[5]_net_1\, Y => \ByteDout_RNO_7[2]_net_1\);
    
    \ByteDout_RNO_0[7]\ : NOR3B
      port map(A => \ByteDout_RNO_3[7]_net_1\, B => 
        \ByteDout_8_i_0[7]\, C => N_708, Y => \ByteDout_8_i_2[7]\);
    
    \CRC_Reg_RNO[9]\ : NOR3
      port map(A => N_440, B => \CRC_Reg_14_i_0_0[9]\, C => N_682, 
        Y => \CRC_Reg_RNO[9]_net_1\);
    
    \Prstate_RNO[1]\ : NOR3A
      port map(A => CMOS_DrvX_0_LVDSen_1, B => N_1015, C => 
        N_1126, Y => \Prstate_RNO[1]_net_1\);
    
    \CRC_Reg[16]\ : DFN1C0
      port map(D => N_288, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \CRC_Reg[16]_net_1\);
    
    \rowcnt_RNI6SI31[6]\ : OR3B
      port map(A => \rowcnt[5]_net_1\, B => \rowcnt[6]_net_1\, C
         => N_312, Y => N_322);
    
    \CRC_Reg_RNO_2[23]\ : NOR2
      port map(A => N_291, B => \CRC_Reg[23]_net_1\, Y => N_641);
    
    \ByteDout_RNO_2[1]\ : NOR3C
      port map(A => N_1047, B => \ByteDout_RNO_7[1]_net_1\, C => 
        N_1046, Y => \ByteDout_8_i_5[1]\);
    
    \Prstate_RNIN2M8_0[0]\ : OR2B
      port map(A => \Prstate[0]_net_1\, B => \ClkEn_0\, Y => 
        N_329);
    
    \Din_Delay3[1]\ : DFN1E1C0
      port map(D => \Din_Delay2[1]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => \ClkEn_2\, Q => \Din_Delay3[1]_net_1\);
    
    \CRC_Reg_RNO_2[20]\ : NOR2
      port map(A => N_291_0, B => \CRC_Reg[20]_net_1\, Y => N_597);
    
    \rowcnt[4]\ : DFN1E0C0
      port map(D => \rowcnt_RNO[4]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => N_329, Q => \rowcnt[4]_net_1\);
    
    StepCnt_n2_0_i_0_RNO : OR2
      port map(A => N_358, B => N_570, Y => StepCnt_n2_0_i_0_0);
    
    \CRC_Reg[34]\ : DFN1C0
      port map(D => N_29, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \CRC_Reg[34]_net_1\);
    
    \DataClkCnt_RNIN6B6[1]\ : NOR2B
      port map(A => \DataClkCnt[1]_net_1\, B => 
        \DataClkCnt[0]_net_1\, Y => N_298);
    
    \CRC_Reg[39]\ : DFN1C0
      port map(D => N_234, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \CRC_Reg[39]_net_1\);
    
    \CRC_Reg[1]\ : DFN1C0
      port map(D => \CRC_Reg_RNO[1]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \CRC_Reg[1]_net_1\);
    
    \DelayCnt_RNO[0]\ : AXOI4
      port map(A => un1_Prstate_3_i, B => \ClkEn_1\, C => 
        DelayCnt_c0, Y => N_146);
    
    \ByteSel_RNITH77[1]\ : NOR2B
      port map(A => \ByteSel[1]_net_1\, B => \ByteSel[0]_net_1\, 
        Y => data_reg30);
    
    \rowcnt_RNO[4]\ : AX1C
      port map(A => N_304, B => \rowcnt[3]_net_1\, C => 
        \rowcnt[4]_net_1\, Y => \rowcnt_RNO[4]_net_1\);
    
    \ByteDout_RNO[6]\ : NOR3C
      port map(A => \ByteDout_RNO_0[6]_net_1\, B => 
        \ByteDout_RNO_1[6]_net_1\, C => \ByteDout_8_i_4[6]\, Y
         => N_184_i_0);
    
    \Shifter_RNO[7]\ : MX2
      port map(A => \Shifter[8]_net_1\, B => \TenbitDout[7]\, S
         => \PtS_En\, Y => \Shifter_4[7]\);
    
    \Prstate[4]\ : DFN1C0
      port map(D => \Prstate_ns[3]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \Prstate[4]_net_1\);
    
    \Shifter_RNO[8]\ : MX2
      port map(A => \Shifter[9]_net_1\, B => \TenbitDout[8]\, S
         => \PtS_En\, Y => \Shifter_4[8]\);
    
    \DataClkCnt_RNO[9]\ : OR3C
      port map(A => N_997, B => N_998, C => N_999, Y => 
        DataClkCnt_e9);
    
    \ByteDout[3]\ : DFN1E1P0
      port map(D => N_178_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        PRE => PLL_Test1_0_SysRst_O, E => N_721, Q => 
        \ByteDout[3]_net_1\);
    
    \ByteSel[0]\ : DFN1C0
      port map(D => ByteSel_n0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \ByteSel[0]_net_1\);
    
    \CRC_Reg_RNO_0[38]\ : AO1D
      port map(A => N_692_0, B => \CRC_Reg[30]_net_1\, C => 
        \CRC_Reg_14_2_i_0[38]\, Y => \CRC_Reg_14_2_i_1[38]\);
    
    \CRC_Reg_RNO_2[31]\ : NOR2
      port map(A => N_291_0, B => \CRC_Reg[31]_net_1\, Y => N_593);
    
    \PKGCnt[2]\ : DFN1E0C0
      port map(D => \PKGCnt_RNO[2]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => N_329_0, Q => \PKGCnt[2]_net_1\);
    
    \DataClkCnt_RNO[1]\ : NOR2B
      port map(A => DataClkCnt_e1_i_0_0, B => N_979, Y => 
        N_16_i_0);
    
    \CRC_Reg_RNO_1[6]\ : NOR2
      port map(A => N_448, B => \CRC_Reg[6]_net_1\, Y => N_607);
    
    \FrameCnt_RNO[5]\ : XOR2
      port map(A => N_327, B => \FrameCnt[5]_net_1\, Y => 
        \FrameCnt_RNO[5]_net_1\);
    
    \ByteDout_RNO_10[2]\ : AO1A
      port map(A => \DelayCnt[2]_net_1\, B => \PKGCnt[13]_net_1\, 
        C => \DelayCnt[1]_net_1\, Y => \ByteDout_8_i_0_a5_0[2]\);
    
    \PKGCnt_RNO[14]\ : AX1
      port map(A => N_347, B => \PKGCnt[13]_net_1\, C => 
        \PKGCnt[14]_net_1\, Y => PKGCnt_n14);
    
    \CRC_Reg_RNO_2[8]\ : NOR2
      port map(A => N_291, B => \CRC_Reg[8]_net_1\, Y => N_629);
    
    \ByteDout_RNO_0[2]\ : NOR3C
      port map(A => N_633, B => \ByteDout_RNO_4[2]_net_1\, C => 
        \ByteDout_RNO_5[2]_net_1\, Y => \ByteDout_8_i_0_1[2]\);
    
    \Prstate_RNO_2[4]\ : NOR2B
      port map(A => \Prstate[5]_net_1\, B => \DelayCnt[3]_net_1\, 
        Y => \Prstate_ns_0_a5_0_0[3]\);
    
    \DataClkCnt_RNO_1[7]\ : NOR2A
      port map(A => \ClkEn_1\, B => N_323, Y => N_992);
    
    \rowcnt[7]\ : DFN1E0C0
      port map(D => N_444_i_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => N_329, Q => 
        \rowcnt[7]_net_1\);
    
    \DataClkCnt_RNO[10]\ : AO1B
      port map(A => N_363, B => \DataClkCnt[10]_net_1\, C => 
        N_1001, Y => DataClkCnt_e10);
    
    \ByteDout_RNO_5[0]\ : OR3A
      port map(A => \ByteDout_8_1_a5_3_0[0]\, B => N_691, C => 
        N_696, Y => N_1037);
    
    \DelayCnt_RNIRIT9[0]\ : OR2B
      port map(A => DelayCnt_c0, B => \ClkEn_1\, Y => N_356);
    
    \ByteDout_RNO_5[7]\ : NOR2
      port map(A => \PKGCnt[2]_net_1\, B => \DelayCnt[2]_net_1\, 
        Y => \ByteDout_8_i_a5_0_0[7]\);
    
    \ByteDout_RNO_2[5]\ : OA1
      port map(A => \FrameCnt[1]_net_1\, B => N_709, C => 
        \ByteDout_RNO_5[5]_net_1\, Y => \ByteDout_8_i_2[5]\);
    
    \rowcnt_RNI26HV1[10]\ : OR2
      port map(A => N_362, B => N_329_0, Y => N_365);
    
    \ByteDout_RNO_4[5]\ : OR2A
      port map(A => \Prstate[4]_net_1\, B => \Fifo_dout[5]\, Y
         => \ByteDout_RNO_4[5]_net_1\);
    
    LVDS_O : DFN1C0
      port map(D => \Shifter[0]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => LVDS_O_c);
    
    \PKGCnt[8]\ : DFN1E0C0
      port map(D => N_449_i_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => N_329, Q => 
        \PKGCnt[8]_net_1\);
    
    \data_reg[6]\ : DFN1C0
      port map(D => data_reg28, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \data_reg[6]_net_1\);
    
    \CRC_Reg[26]\ : DFN1C0
      port map(D => \CRC_Reg_RNO[26]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \CRC_Reg[26]_net_1\);
    
    tok : DFN1E1C0
      port map(D => N_746, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => \ClkEn\, Q => tok_c);
    
    \CRC_Reg_RNO[25]\ : OA1B
      port map(A => \CRC_Reg[25]_net_1\, B => N_291_0, C => 
        \CRC_Reg_14_i_0_1[25]\, Y => N_17);
    
    \rowcnt_RNO[3]\ : XOR2
      port map(A => \rowcnt[3]_net_1\, B => N_304, Y => 
        \rowcnt_RNO[3]_net_1\);
    
    \FrameCnt_RNIMCLA[4]\ : NOR3C
      port map(A => \FrameCnt[3]_net_1\, B => N_320, C => 
        \FrameCnt[4]_net_1\, Y => N_327);
    
    \PKGCnt_RNO[5]\ : XOR2
      port map(A => \PKGCnt[5]_net_1\, B => N_300, Y => 
        \PKGCnt_RNO[5]_net_1\);
    
    \CRC_Reg_RNO[17]\ : NOR3
      port map(A => \CRC_Reg_14_i_0_0[17]\, B => N_674, C => 
        N_673, Y => \CRC_Reg_RNO[17]_net_1\);
    
    \CRC_Reg_RNO[8]\ : NOR3
      port map(A => N_436, B => \CRC_Reg_14_2_i_0[8]\, C => N_629, 
        Y => N_256);
    
    \ByteDout_RNO_1[7]\ : OR2
      port map(A => \rowcnt[7]_net_1\, B => N_705, Y => 
        \ByteDout_RNO_1[7]_net_1\);
    
    \Shifter_RNO[1]\ : MX2
      port map(A => \Shifter[2]_net_1\, B => \TenbitDout[1]\, S
         => \PtS_En\, Y => \Shifter_4[1]\);
    
    \Din_Delay2[4]\ : DFN1E1P0
      port map(D => \Din_Delay1[4]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, PRE => PLL_Test1_0_SysRst_O, E
         => \ClkEn_2\, Q => \Din_Delay2[4]_net_1\);
    
    \DataClkCnt_RNO[6]\ : NOR2A
      port map(A => N_979, B => DataClkCnt_e6_i_0_0, Y => N_26);
    
    \ByteDout[2]\ : DFN1E1P0
      port map(D => N_12_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, PRE
         => PLL_Test1_0_SysRst_O, E => N_721, Q => 
        \ByteDout[2]_net_1\);
    
    \Din_Delay2[5]\ : DFN1E1P0
      port map(D => \Din_Delay1[5]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, PRE => PLL_Test1_0_SysRst_O, E
         => \ClkEn_2\, Q => \Din_Delay2[5]_net_1\);
    
    \CRC_Reg_RNO[2]\ : OA1B
      port map(A => \CRC_Reg[2]_net_1\, B => N_448, C => 
        \CRC_Reg_14_i_0_1[2]\, Y => \CRC_Reg_RNO[2]_net_1\);
    
    \CRC_Reg_RNO_0[18]\ : XA1A
      port map(A => \CRC_Reg[39]_net_1\, B => \CRC_Reg[17]_net_1\, 
        C => N_690, Y => N_438);
    
    \StepCnt_RNI3G91[1]\ : NOR2B
      port map(A => \StepCnt[1]_net_1\, B => \StepCnt[0]_net_1\, 
        Y => N_341);
    
    \Din_Delay3[4]\ : DFN1E1P0
      port map(D => \Din_Delay2[4]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, PRE => PLL_Test1_0_SysRst_O, E
         => \ClkEn_2\, Q => \Din_Delay3[4]_net_1\);
    
    \Din_Delay3[6]\ : DFN1E1C0
      port map(D => \Din_Delay2[6]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => \ClkEn\, Q => \Din_Delay3[6]_net_1\);
    
    \FrameCnt[2]\ : DFN1E0C0
      port map(D => \FrameCnt_RNO[2]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => N_365, Q => \FrameCnt[2]_net_1\);
    
    \CRC_Reg_RNO_1[39]\ : AO1C
      port map(A => \CRC_Reg[38]_net_1\, B => N_690_0, C => 
        CMOS_DrvX_0_LVDSen_0, Y => \CRC_Reg_14_2_i_0[39]\);
    
    CRC_ResultAva_RNO_3 : NOR3A
      port map(A => \Prstate[1]_net_1\, B => \DelayCnt[2]_net_1\, 
        C => \DelayCnt[3]_net_1\, Y => CRC_ResultAva_3_0_o2_0);
    
    StepCnt_n2_0_i_0_a5 : NOR2
      port map(A => N_341, B => \StepCnt[2]_net_1\, Y => N_570);
    
    \FrameCnt_RNO[0]\ : XNOR2
      port map(A => \FrameCnt[0]_net_1\, B => N_365, Y => 
        \FrameCnt_RNO[0]_net_1\);
    
    \ClkDivCnt_RNILBNB[1]\ : OR2A
      port map(A => \ClkDivCnt[0]_net_1\, B => 
        \ClkDivCnt[1]_net_1\, Y => bit_en2_1);
    
    \CRC_Reg_RNO[36]\ : OA1B
      port map(A => \CRC_Reg[36]_net_1\, B => N_291_0, C => 
        \CRC_Reg_14_i_0_1[36]\, Y => N_33);
    
    \ByteDout_RNO_5[4]\ : OR2A
      port map(A => \Prstate[4]_net_1\, B => \Fifo_dout[4]\, Y
         => \ByteDout_RNO_5[4]_net_1\);
    
    \PKGCnt_RNIT2SE1[8]\ : NOR2A
      port map(A => \PKGCnt[8]_net_1\, B => N_310, Y => N_316);
    
    \CRC_Reg_RNO_1[25]\ : AO1C
      port map(A => \CRC_Reg[24]_net_1\, B => N_690_0, C => 
        CMOS_DrvX_0_LVDSen_1, Y => \CRC_Reg_14_i_0_0[25]\);
    
    \ClkDivCnt_RNO[1]\ : OA1A
      port map(A => clkdivcnt7_0, B => bit_en2_1, C => I_5, Y => 
        \ClkDivCnt_3[1]\);
    
    \CRC_Reg_RNO_1[27]\ : NOR2
      port map(A => N_692, B => \CRC_Reg[19]_net_1\, Y => N_659);
    
    \CRC_Reg[3]\ : DFN1C0
      port map(D => \CRC_Reg_RNO[3]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \CRC_Reg[3]_net_1\);
    
    \CRC_Reg_RNO_1[26]\ : NOR2
      port map(A => N_692, B => \CRC_Reg[18]_net_1\, Y => N_662);
    
    \ByteDout_RNO[3]\ : NOR3C
      port map(A => \ByteDout_RNO_0[3]_net_1\, B => 
        \ByteDout_8_i_1[3]\, C => \ByteDout_RNO_2[3]_net_1\, Y
         => N_178_i_0);
    
    \rowcnt[1]\ : DFN1E0C0
      port map(D => N_385_i, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => N_329, Q => 
        \rowcnt[1]_net_1\);
    
    \CRC_Reg_RNO_2[18]\ : NOR2
      port map(A => N_291, B => \CRC_Reg[18]_net_1\, Y => N_670);
    
    \Prstate[0]\ : DFN1C0
      port map(D => \Prstate_ns[7]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \Prstate[0]_net_1\);
    
    \Din_Delay3[0]\ : DFN1E1C0
      port map(D => \Din_Delay2[0]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => \ClkEn_2\, Q => \Din_Delay3[0]_net_1\);
    
    \data_reg[0]\ : DFN1C0
      port map(D => data_reg27, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \data_reg[0]_net_1\);
    
    REen_RNO : AO1
      port map(A => REen_1_0_0_a5_0, B => \REen\, C => 
        \Prstate[5]_net_1\, Y => REen_1);
    
    \Din_Delay3[3]\ : DFN1E1P0
      port map(D => \Din_Delay2[3]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, PRE => PLL_Test1_0_SysRst_O, E
         => \ClkEn_2\, Q => \Din_Delay3[3]_net_1\);
    
    \CRC_Reg_RNO_1[21]\ : AO1C
      port map(A => \CRC_Reg[20]_net_1\, B => N_690_0, C => 
        CMOS_DrvX_0_LVDSen_0, Y => \CRC_Reg_14_2_i_0[21]\);
    
    \CRC_Reg_RNO_1[15]\ : OAI1
      port map(A => \CRC_Reg[7]_net_1\, B => N_692, C => 
        CMOS_DrvX_0_LVDSen_1, Y => \CRC_Reg_14_2_i_0[15]\);
    
    \Prstate_RNO_1[5]\ : NOR3
      port map(A => N_696, B => \Prstate_ns_i_0_0_a5_0_0[2]\, C
         => N_356, Y => N_1014);
    
    \CRC_Reg_RNO_1[17]\ : NOR2
      port map(A => N_692, B => \CRC_Reg[9]_net_1\, Y => N_674);
    
    \CRC_Reg_RNO_0[29]\ : AO1D
      port map(A => N_692_0, B => \CRC_Reg[21]_net_1\, C => 
        \CRC_Reg_14_2_i_0[29]\, Y => \CRC_Reg_14_2_i_1[29]\);
    
    \DataClkCnt_RNO[4]\ : NOR2A
      port map(A => N_979, B => DataClkCnt_e4_i_0_0, Y => N_22);
    
    \Shifter[9]\ : DFN1E1C0
      port map(D => \TenbitDout[9]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => \PtS_En\, Q => \Shifter[9]_net_1\);
    
    \CRC_Reg[30]\ : DFN1C0
      port map(D => N_238, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \CRC_Reg[30]_net_1\);
    
    \DataClkCnt_RNIHK1J[5]\ : NOR2B
      port map(A => N_309, B => \DataClkCnt[5]_net_1\, Y => N_314);
    
    \CRC_Reg_RNO_1[16]\ : OAI1
      port map(A => \CRC_Reg[8]_net_1\, B => N_692, C => 
        CMOS_DrvX_0_LVDSen_1, Y => \CRC_Reg_14_2_i_0[16]\);
    
    \Prstate_RNO_1[4]\ : OR3B
      port map(A => CMOS_DrvX_0_LVDSen_1, B => \Prstate[4]_net_1\, 
        C => N_355, Y => N_1082);
    
    \Shifter_RNO[2]\ : MX2
      port map(A => \Shifter[3]_net_1\, B => \TenbitDout[2]\, S
         => \PtS_En\, Y => \Shifter_4[2]\);
    
    \CRC_Reg_RNO_1[0]\ : NOR2A
      port map(A => N_450, B => \CRC_Reg[0]_net_1\, Y => N_576);
    
    \PKGCnt_RNO[8]\ : XNOR2
      port map(A => \PKGCnt[8]_net_1\, B => N_310, Y => 
        N_449_i_i_0);
    
    \CRC_Reg[0]\ : DFN1C0
      port map(D => \CRC_Reg_RNO[0]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \CRC_Reg[0]_net_1\);
    
    \ByteDout_RNO[4]\ : NOR3C
      port map(A => \ByteDout_8_i_2[4]\, B => 
        \ByteDout_RNO_1[4]_net_1\, C => \ByteDout_8_i_3[4]\, Y
         => N_180_i_0);
    
    \CRC_Reg[8]\ : DFN1C0
      port map(D => N_256, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \CRC_Reg[8]_net_1\);
    
    \ByteDout_RNO_5[6]\ : OR3
      port map(A => \Prstate[4]_net_1\, B => \Prstate[5]_net_1\, 
        C => N_368, Y => N_1067);
    
    \Prstate_RNO[0]\ : OA1
      port map(A => N_1126, B => \Prstate_RNO_0[0]_net_1\, C => 
        CMOS_DrvX_0_LVDSen_2, Y => \Prstate_ns[7]\);
    
    \CRC_Reg[15]\ : DFN1C0
      port map(D => N_290, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \CRC_Reg[15]_net_1\);
    
    \ByteDout_RNO[5]\ : NOR3C
      port map(A => \ByteDout_RNO_0[5]_net_1\, B => 
        \ByteDout_8_i_1[5]\, C => \ByteDout_8_i_2[5]\, Y => 
        N_182_i_0);
    
    \Prstate[1]\ : DFN1C0
      port map(D => \Prstate_RNO[1]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \Prstate[1]_net_1\);
    
    \CRC_Reg[7]\ : DFN1C0
      port map(D => \CRC_Reg_RNO[7]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \CRC_Reg[7]_net_1\);
    
    \StepCnt_RNIA7K6[3]\ : NOR2
      port map(A => \StepCnt[3]_net_1\, B => \ClkEn_0\, Y => 
        N_690_0);
    
    Com_8b10b : enc_8b10b
      port map(TenbitDout(9) => \TenbitDout[9]\, TenbitDout(8)
         => \TenbitDout[8]\, TenbitDout(7) => \TenbitDout[7]\, 
        TenbitDout(6) => \TenbitDout[6]\, TenbitDout(5) => 
        \TenbitDout[5]\, TenbitDout(4) => \TenbitDout[4]\, 
        TenbitDout(3) => \TenbitDout[3]\, TenbitDout(2) => 
        \TenbitDout[2]\, TenbitDout(1) => \TenbitDout[1]\, 
        TenbitDout(0) => \TenbitDout[0]\, Din_Delay4_6 => 
        \Din_Delay4[6]_net_1\, Din_Delay4_5 => 
        \Din_Delay4[5]_net_1\, Din_Delay4_7 => 
        \Din_Delay4[7]_net_1\, Din_Delay4_2 => 
        \Din_Delay4[2]_net_1\, Din_Delay4_0 => 
        \Din_Delay4[0]_net_1\, Din_Delay4_1 => 
        \Din_Delay4[1]_net_1\, CRC_Reg_6 => \CRC_Reg[38]_net_1\, 
        CRC_Reg_5 => \CRC_Reg[37]_net_1\, CRC_Reg_7 => 
        \CRC_Reg[39]_net_1\, CRC_Reg_2 => \CRC_Reg[34]_net_1\, 
        CRC_Reg_0 => \CRC_Reg[32]_net_1\, CRC_Reg_1 => 
        \CRC_Reg[33]_net_1\, Bit_En => \Bit_En\, 
        PLL_Test1_0_SysRst_O => PLL_Test1_0_SysRst_O, 
        PLL_Test1_0_Sys_66M_Clk => PLL_Test1_0_Sys_66M_Clk, 
        Kin_Delay4 => \Kin_Delay4\, CRC_ResultAva => 
        \CRC_ResultAva\, N_423 => N_423, N_422 => N_422, N_425
         => N_425, N_426 => N_426);
    
    \ClkDivCnt[3]\ : DFN1C0
      port map(D => \ClkDivCnt_3[3]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \ClkDivCnt[3]_net_1\);
    
    \FrameCnt_RNO[3]\ : XOR2
      port map(A => N_320, B => \FrameCnt[3]_net_1\, Y => 
        \FrameCnt_RNO[3]_net_1\);
    
    \DataClkCnt_RNO[0]\ : AXOI5
      port map(A => N_5, B => \ClkEn_1\, C => 
        \DataClkCnt[0]_net_1\, Y => N_7_0);
    
    \PKGCnt_RNIM0KF[2]\ : OR3C
      port map(A => \PKGCnt[0]_net_1\, B => \PKGCnt[1]_net_1\, C
         => \PKGCnt[2]_net_1\, Y => N_295);
    
    ClkEn_1_RNIF8SQ : OR3B
      port map(A => CMOS_DrvX_0_LVDSen_2, B => N_450, C => N_690, 
        Y => StepCnte);
    
    \CRC_Reg_RNO_1[11]\ : NOR2
      port map(A => N_692, B => \CRC_Reg[3]_net_1\, Y => N_677);
    
    \CRC_Reg_RNO_1[22]\ : NOR2
      port map(A => N_692, B => \CRC_Reg[14]_net_1\, Y => N_639);
    
    \DelayCnt_RNI1M8L_0[2]\ : OR3
      port map(A => N_313, B => N_693, C => \DelayCnt[2]_net_1\, 
        Y => N_709);
    
    \Shifter[3]\ : DFN1C0
      port map(D => \Shifter_4[3]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \Shifter[3]_net_1\);
    
    \Prstate_RNO_0[2]\ : NOR2B
      port map(A => \Prstate[2]_net_1\, B => CMOS_DrvX_0_LVDSen_1, 
        Y => \Prstate_ns_0_a5_0[5]\);
    
    \CRC_Reg[6]\ : DFN1C0
      port map(D => \CRC_Reg_RNO[6]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \CRC_Reg[6]_net_1\);
    
    \ByteDout_RNO_0[3]\ : OR3
      port map(A => DelayCnt_c0, B => N_693, C => N_414, Y => 
        \ByteDout_RNO_0[3]_net_1\);
    
    \StepCnt_RNO_0[3]\ : XOR2
      port map(A => \StepCnt[3]_net_1\, B => N_358, Y => 
        N_394_i_i_0);
    
    \DataClkCnt[3]\ : DFN1C0
      port map(D => N_20, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \DataClkCnt[3]_net_1\);
    
    \CRC_Reg_RNO_0[1]\ : OR3
      port map(A => N_623, B => N_624, C => N_353, Y => 
        \CRC_Reg_14_i_0_1[1]\);
    
    \CRC_Reg_RNO[35]\ : OA1B
      port map(A => \CRC_Reg[35]_net_1\, B => N_291_0, C => 
        \CRC_Reg_14_i_0_1[35]\, Y => N_31);
    
    \FrameCnt_RNINQC6[2]\ : NOR3C
      port map(A => \FrameCnt[0]_net_1\, B => \FrameCnt[1]_net_1\, 
        C => \FrameCnt[2]_net_1\, Y => N_320);
    
    \CRC_Reg_RNO_2[34]\ : NOR2
      port map(A => N_291, B => \CRC_Reg[34]_net_1\, Y => N_650);
    
    \ByteDout_RNO_4[4]\ : OR3
      port map(A => N_704, B => \FrameCnt[8]_net_1\, C => N_698, 
        Y => \ByteDout_RNO_4[4]_net_1\);
    
    ClkEn_1_RNI218K : NAND2
      port map(A => CMOS_DrvX_0_LVDSen_0, B => N_450, Y => 
        un1_StepCnt_3_i_0);
    
    \ByteDout_RNO_10[1]\ : NOR2A
      port map(A => \FrameCnt[5]_net_1\, B => DelayCnt_c0, Y => 
        N_376);
    
    Kin : DFN1E1P0
      port map(D => N_970, CLK => PLL_Test1_0_Sys_66M_Clk, PRE
         => PLL_Test1_0_SysRst_O, E => \ClkEn\, Q => \Kin\);
    
    \ByteDout_RNO_6[3]\ : MX2
      port map(A => \PKGCnt[14]_net_1\, B => \FrameCnt[7]_net_1\, 
        S => \DelayCnt[1]_net_1\, Y => N_413);
    
    \PKGCnt_RNO[11]\ : XOR2
      port map(A => N_325, B => \PKGCnt[11]_net_1\, Y => 
        PKGCnt_n11);
    
    LVDS_ok_RNIGAO5 : INV
      port map(A => \FrameMk_0_LVDS_ok\, Y => FrameMk_0_LVDS_ok_i);
    
    CRC_ResultAva_RNO_0 : NOR3B
      port map(A => \Prstate[2]_net_1\, B => \DelayCnt[2]_net_1\, 
        C => DelayCnt_c0, Y => CRC_ResultAva_3_0_a5_0_2);
    
    \ByteDout_RNO[1]\ : NOR3C
      port map(A => N_1045, B => \ByteDout_8_i_2[1]\, C => 
        \ByteDout_8_i_5[1]\, Y => N_176_i_0);
    
    un1_clkdivcnt_I_9 : XOR2
      port map(A => N_7, B => \ClkDivCnt[2]_net_1\, Y => I_9);
    
    \DataClkCnt_RNO_3[11]\ : NOR2A
      port map(A => \DataClkCnt[11]_net_1\, B => 
        \DataClkCnt[10]_net_1\, Y => DataClkCnt_e11_0_0_a5_0_0);
    
    \DelayCnt_RNO[3]\ : NOR2
      port map(A => N_1019, B => N_398_i, Y => N_188);
    
    \CRC_Reg_RNO_1[12]\ : OAI1
      port map(A => \CRC_Reg[4]_net_1\, B => N_692_0, C => 
        CMOS_DrvX_0_LVDSen_0, Y => \CRC_Reg_14_2_i_0[12]\);
    
    \PKGCnt_RNO[2]\ : AX1C
      port map(A => \PKGCnt[0]_net_1\, B => \PKGCnt[1]_net_1\, C
         => \PKGCnt[2]_net_1\, Y => \PKGCnt_RNO[2]_net_1\);
    
    \CRC_Reg[25]\ : DFN1C0
      port map(D => N_17, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \CRC_Reg[25]_net_1\);
    
    \CRC_Reg_RNO[24]\ : NOR3
      port map(A => N_441, B => \CRC_Reg_14_2_i_0[24]\, C => 
        N_684, Y => N_286);
    
    \ByteDout_RNO_7[0]\ : OR2B
      port map(A => \Prstate[4]_net_1\, B => \Fifo_dout[0]\, Y
         => N_1035);
    
    \ByteDout_RNO_6[0]\ : OR3A
      port map(A => N_368, B => \Prstate[4]_net_1\, C => 
        \Prstate[5]_net_1\, Y => N_1034);
    
    \CRC_Reg_RNO_2[2]\ : NOR2A
      port map(A => N_690, B => \CRC_Reg[1]_net_1\, Y => N_621);
    
    \ByteDout_RNO_8[0]\ : MX2
      port map(A => \FrameCnt[4]_net_1\, B => \rowcnt[8]_net_1\, 
        S => \DelayCnt[2]_net_1\, Y => N_412);
    
    \ClkDivCnt_RNIPRNB[3]\ : NOR2A
      port map(A => \ClkDivCnt[3]_net_1\, B => 
        \ClkDivCnt[2]_net_1\, Y => clkdivcnt7_0);
    
    \ByteDout_RNO_5[5]\ : OR2
      port map(A => \rowcnt[5]_net_1\, B => N_705, Y => 
        \ByteDout_RNO_5[5]_net_1\);
    
    \CRC_Reg_RNO_2[6]\ : NOR2A
      port map(A => N_690_0, B => \CRC_Reg[5]_net_1\, Y => N_609);
    
    \CRC_Reg_RNO_2[30]\ : NOR2
      port map(A => N_291_0, B => \CRC_Reg[30]_net_1\, Y => N_595);
    
    WE : DFN1C0
      port map(D => Main_ctl4SD_0_ByteRdEn, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \WE\);
    
    CRC_ResultAva_RNIS5FH : OR2A
      port map(A => N_692, B => N_690, Y => N_291);
    
    \DataClkCnt_RNIIDMC[3]\ : NOR2B
      port map(A => N_302, B => \DataClkCnt[3]_net_1\, Y => N_305);
    
    \PKGCnt[9]\ : DFN1E0C0
      port map(D => PKGCnt_n9, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => N_329, Q => 
        \PKGCnt[9]_net_1\);
    
    \ByteDout_RNO_11[1]\ : OR2
      port map(A => \rowcnt[1]_net_1\, B => N_313, Y => 
        \ByteDout_8_i_a5_4_0[1]\);
    
    Kin_Delay3 : DFN1E1P0
      port map(D => \Kin_Delay2\, CLK => PLL_Test1_0_Sys_66M_Clk, 
        PRE => PLL_Test1_0_SysRst_O, E => \ClkEn\, Q => 
        \Kin_Delay3\);
    
    \ClkDivCnt_RNO[3]\ : OA1A
      port map(A => clkdivcnt7_0, B => bit_en2_1, C => I_13, Y
         => \ClkDivCnt_3[3]\);
    
    \FrameCnt[0]\ : DFN1C0
      port map(D => \FrameCnt_RNO[0]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \FrameCnt[0]_net_1\);
    
    \ByteDout_RNO_5[2]\ : OR3
      port map(A => DelayCnt_c0, B => N_693, C => 
        \ByteDout_8_i_0_a5_2_0[2]\, Y => 
        \ByteDout_RNO_5[2]_net_1\);
    
    \rowcnt_RNO[7]\ : XNOR2
      port map(A => \rowcnt[7]_net_1\, B => N_322, Y => 
        N_444_i_i_0);
    
    \DelayCnt_RNIBRS7[1]\ : OR2A
      port map(A => \DelayCnt[1]_net_1\, B => \DelayCnt[2]_net_1\, 
        Y => N_704);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    \DelayCnt_RNO_0[1]\ : NOR2A
      port map(A => N_356, B => \DelayCnt[1]_net_1\, Y => N_1017);
    
    \DataClkCnt[9]\ : DFN1C0
      port map(D => DataClkCnt_e9, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \DataClkCnt[9]_net_1\);
    
    \rowcnt_RNO[9]\ : XNOR2
      port map(A => N_334, B => \rowcnt[9]_net_1\, Y => rowcnt_n9);
    
    \DataClkCnt_RNI287M[6]\ : NOR2B
      port map(A => N_314, B => \DataClkCnt[6]_net_1\, Y => N_318);
    
    \DataClkCnt_RNI9UM81[3]\ : NOR3C
      port map(A => DataOk_0_sqmuxa_0_a2_0_a5_8, B => 
        DataOk_0_sqmuxa_0_a2_0_a5_7, C => 
        DataOk_0_sqmuxa_0_a2_0_a5_9, Y => DataOk_0_sqmuxa);
    
    \DelayCnt_RNI2DD9_0[3]\ : OR2
      port map(A => N_691, B => \DelayCnt[3]_net_1\, Y => N_693);
    
    \CRC_Reg_RNO_1[35]\ : AO1C
      port map(A => \CRC_Reg[34]_net_1\, B => N_690_0, C => 
        CMOS_DrvX_0_LVDSen_0, Y => \CRC_Reg_14_i_0_0[35]\);
    
    \CRC_Reg_RNO[16]\ : NOR3
      port map(A => N_442, B => \CRC_Reg_14_2_i_0[16]\, C => 
        N_686, Y => N_288);
    
    \CRC_Reg_RNO_1[37]\ : AO1C
      port map(A => \CRC_Reg[36]_net_1\, B => N_690_0, C => 
        CMOS_DrvX_0_LVDSen_0, Y => \CRC_Reg_14_2_i_0[37]\);
    
    \ByteDout_RNO_1[2]\ : OR3
      port map(A => DelayCnt_c0, B => N_693, C => N_2220_tz, Y
         => \ByteDout_RNO_1[2]_net_1\);
    
    \StepCnt_RNIB7K6[3]\ : NOR2
      port map(A => \StepCnt[3]_net_1\, B => \ClkEn_1\, Y => 
        N_690);
    
    \CRC_Reg_RNO_1[36]\ : AO1C
      port map(A => \CRC_Reg[35]_net_1\, B => N_690_0, C => 
        CMOS_DrvX_0_LVDSen_0, Y => \CRC_Reg_14_i_0_0[36]\);
    
    \PKGCnt_RNI0M012[12]\ : OR3C
      port map(A => N_325, B => \PKGCnt[11]_net_1\, C => 
        \PKGCnt[12]_net_1\, Y => N_347);
    
    \Din_Delay1[1]\ : DFN1E1C0
      port map(D => \ByteDout[1]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => \ClkEn_1\, Q => \Din_Delay1[1]_net_1\);
    
    \PKGCnt_RNIPJCO1[10]\ : NOR3C
      port map(A => N_316, B => \PKGCnt[9]_net_1\, C => 
        \PKGCnt[10]_net_1\, Y => N_325);
    
    un1_clkdivcnt_I_12 : AND3
      port map(A => \ClkDivCnt[0]_net_1\, B => 
        \ClkDivCnt[1]_net_1\, C => \ClkDivCnt[2]_net_1\, Y => N_4);
    
    \PKGCnt_RNICNE41[6]\ : NOR3C
      port map(A => N_300, B => \PKGCnt[5]_net_1\, C => 
        \PKGCnt[6]_net_1\, Y => N_306);
    
    \ByteDout_RNO_6[4]\ : OR2A
      port map(A => N_708, B => \PKGCnt[15]_net_1\, Y => N_1055);
    
    \Din_Delay3[7]\ : DFN1E1P0
      port map(D => \Din_Delay2[7]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, PRE => PLL_Test1_0_SysRst_O, E
         => \ClkEn\, Q => \Din_Delay3[7]_net_1\);
    
    \DataClkCnt_RNO_2[11]\ : OR2B
      port map(A => DataClkCnt_e11_0_0_a5_0_0, B => N_5, Y => 
        N_1004);
    
    \ByteDout_RNO_3[6]\ : NOR3C
      port map(A => N_1067, B => \ByteDout_RNO_6[6]_net_1\, C => 
        N_1068, Y => \ByteDout_8_i_1[6]\);
    
    \DataClkCnt[1]\ : DFN1C0
      port map(D => N_16_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \DataClkCnt[1]_net_1\);
    
    \DataClkCnt_RNO_2[8]\ : OR3
      port map(A => N_706_i, B => \DataClkCnt[8]_net_1\, C => 
        N_323, Y => N_995);
    
    \rowcnt[2]\ : DFN1E0C0
      port map(D => N_392_i_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => N_329, Q => 
        \rowcnt[2]_net_1\);
    
    \Prstate_RNO[4]\ : AO1C
      port map(A => N_356, B => \Prstate_ns_0_a5_0_2[3]\, C => 
        N_1082, Y => \Prstate_ns[3]\);
    
    \CRC_Reg_RNO_1[24]\ : OAI1
      port map(A => \CRC_Reg[16]_net_1\, B => N_692, C => 
        CMOS_DrvX_0_LVDSen_1, Y => \CRC_Reg_14_2_i_0[24]\);
    
    \ByteDout[1]\ : DFN1E1C0
      port map(D => N_176_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => N_721, Q => 
        \ByteDout[1]_net_1\);
    
    \CRC_Reg_RNO_1[31]\ : OAI1
      port map(A => \CRC_Reg[23]_net_1\, B => N_692_0, C => 
        CMOS_DrvX_0_LVDSen_0, Y => \CRC_Reg_14_2_i_0[31]\);
    
    \rowcnt_RNO[2]\ : AX1C
      port map(A => \rowcnt[0]_net_1\, B => \rowcnt[1]_net_1\, C
         => \rowcnt[2]_net_1\, Y => N_392_i_i_0);
    
    CRC_ResultAva : DFN1E1C0
      port map(D => CRC_ResultAva_3, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => \ClkEn_1\, Q => \CRC_ResultAva\);
    
    \CRC_Reg[18]\ : DFN1C0
      port map(D => \CRC_Reg_RNO[18]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \CRC_Reg[18]_net_1\);
    
    un1_clkdivcnt_I_5 : XOR2
      port map(A => \ClkDivCnt[0]_net_1\, B => 
        \ClkDivCnt[1]_net_1\, Y => I_5);
    
    \ByteDout[5]\ : DFN1E1P0
      port map(D => N_182_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        PRE => PLL_Test1_0_SysRst_O, E => N_721, Q => 
        \ByteDout[5]_net_1\);
    
    \CRC_Reg_RNO_0[5]\ : AO1D
      port map(A => N_450, B => \ByteDout[5]_net_1\, C => N_612, 
        Y => \CRC_Reg_14_i_0_0[5]\);
    
    ClkEn : DFN1C0
      port map(D => clken2, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \ClkEn\);
    
    \CRC_Reg[36]\ : DFN1C0
      port map(D => N_33, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \CRC_Reg[36]_net_1\);
    
    CRC_ResultAva_RNIFHTG : OR2B
      port map(A => N_692, B => CMOS_DrvX_0_LVDSen_2, Y => N_353);
    
    \CRC_Reg_RNO_0[25]\ : AO1D
      port map(A => N_692, B => \CRC_Reg[17]_net_1\, C => 
        \CRC_Reg_14_i_0_0[25]\, Y => \CRC_Reg_14_i_0_1[25]\);
    
    \CRC_Reg_RNO_2[1]\ : NOR2A
      port map(A => N_690, B => \CRC_Reg[0]_net_1\, Y => N_624);
    
    \Shifter_RNO[6]\ : MX2
      port map(A => \Shifter[7]_net_1\, B => \TenbitDout[6]\, S
         => \PtS_En\, Y => \Shifter_4[6]\);
    
    \Din_Delay3[2]\ : DFN1E1P0
      port map(D => \Din_Delay2[2]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, PRE => PLL_Test1_0_SysRst_O, E
         => \ClkEn_2\, Q => \Din_Delay3[2]_net_1\);
    
    \CRC_Reg_RNO_0[27]\ : AO1C
      port map(A => \CRC_Reg[26]_net_1\, B => N_690_0, C => 
        CMOS_DrvX_0_LVDSen_1, Y => \CRC_Reg_14_i_0_0[27]\);
    
    \Din_Delay4[5]\ : DFN1E1P0
      port map(D => \Din_Delay3[5]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, PRE => PLL_Test1_0_SysRst_O, E
         => \ClkEn\, Q => \Din_Delay4[5]_net_1\);
    
    \Din_Delay4[7]\ : DFN1E1P0
      port map(D => \Din_Delay3[7]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, PRE => PLL_Test1_0_SysRst_O, E
         => \ClkEn\, Q => \Din_Delay4[7]_net_1\);
    
    \Din_Delay1[6]\ : DFN1E1C0
      port map(D => \ByteDout[6]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => \ClkEn_2\, Q => \Din_Delay1[6]_net_1\);
    
    \CRC_Reg_RNO[1]\ : OA1B
      port map(A => \CRC_Reg[1]_net_1\, B => N_448, C => 
        \CRC_Reg_14_i_0_1[1]\, Y => \CRC_Reg_RNO[1]_net_1\);
    
    \CRC_Reg_RNO_0[26]\ : AO1C
      port map(A => \CRC_Reg[25]_net_1\, B => N_690_0, C => 
        CMOS_DrvX_0_LVDSen_1, Y => \CRC_Reg_14_i_0_0[26]\);
    
    \CRC_Reg_RNO_1[23]\ : NOR2
      port map(A => N_692, B => \CRC_Reg[15]_net_1\, Y => N_642);
    
    \DataClkCnt_RNO_0[2]\ : AX1E
      port map(A => N_298, B => \ClkEn_0\, C => 
        \DataClkCnt[2]_net_1\, Y => DataClkCnt_e2_i_0_0);
    
    \CRC_Reg_RNO_1[20]\ : OAI1
      port map(A => \CRC_Reg[12]_net_1\, B => N_692_0, C => 
        CMOS_DrvX_0_LVDSen_0, Y => \CRC_Reg_14_2_i_0[20]\);
    
    \ByteDout[0]\ : DFN1E1C0
      port map(D => \ByteDout_8[0]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => N_721, Q => \ByteDout[0]_net_1\);
    
    \DelayCnt[3]\ : DFN1C0
      port map(D => N_188, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \DelayCnt[3]_net_1\);
    
    \CRC_Reg_RNO_1[14]\ : AO1C
      port map(A => \CRC_Reg[13]_net_1\, B => N_690_0, C => 
        CMOS_DrvX_0_LVDSen_0, Y => \CRC_Reg_14_2_i_0[14]\);
    
    \Din_Delay1[2]\ : DFN1E1P0
      port map(D => \ByteDout[2]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, PRE => PLL_Test1_0_SysRst_O, E
         => \ClkEn_1\, Q => \Din_Delay1[2]_net_1\);
    
    Kin_Delay1 : DFN1E1P0
      port map(D => \Kin\, CLK => PLL_Test1_0_Sys_66M_Clk, PRE
         => PLL_Test1_0_SysRst_O, E => \ClkEn\, Q => \Kin_Delay1\);
    
    \CRC_Reg_RNO_1[32]\ : AO1C
      port map(A => \CRC_Reg[31]_net_1\, B => N_690_0, C => 
        CMOS_DrvX_0_LVDSen_0, Y => \CRC_Reg_14_i_0_0[32]\);
    
    Bit_En : DFN1C0
      port map(D => bit_en2, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \Bit_En\);
    
    \DelayCnt_RNO[1]\ : NOR3
      port map(A => N_333_i_0, B => N_1019, C => N_1017, Y => 
        N_148);
    
    \CRC_Reg_RNO_0[21]\ : AO1D
      port map(A => N_692_0, B => \CRC_Reg[13]_net_1\, C => 
        \CRC_Reg_14_2_i_0[21]\, Y => \CRC_Reg_14_2_i_1[21]\);
    
    \ByteDout[4]\ : DFN1E1P0
      port map(D => N_180_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        PRE => PLL_Test1_0_SysRst_O, E => N_721, Q => 
        \ByteDout[4]_net_1\);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    \Din_Delay4[1]\ : DFN1E1C0
      port map(D => \Din_Delay3[1]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => \ClkEn\, Q => \Din_Delay4[1]_net_1\);
    
    \Shifter[1]\ : DFN1C0
      port map(D => \Shifter_4[1]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \Shifter[1]_net_1\);
    
    \Prstate_RNIDOIU[3]\ : OR3C
      port map(A => CMOS_DrvX_0_LVDSen_1, B => 
        \Prstate_ns_0_a5_0_0[5]\, C => N_333_i_0, Y => N_548);
    
    \CRC_Reg_RNO[34]\ : NOR3
      port map(A => N_437, B => \CRC_Reg_14_i_0_0[34]\, C => 
        N_650, Y => N_29);
    
    REen_RNO_0 : NOR2
      port map(A => \Prstate[7]_net_1\, B => \Prstate[3]_net_1\, 
        Y => REen_1_0_0_a5_0);
    
    \ByteDout_RNO_6[2]\ : OA1
      port map(A => \FrameCnt[6]_net_1\, B => N_704, C => 
        \ByteDout_8_i_0_a5_0[2]\, Y => N_2220_tz);
    
    \ByteDout_RNO_3[1]\ : OA1A
      port map(A => \Prstate[4]_net_1\, B => \Fifo_dout[1]\, C
         => N_1042, Y => \ByteDout_8_i_0[1]\);
    
    \ByteDout_RNO_2[3]\ : OR3A
      port map(A => DelayCnt_c0, B => N_702, C => 
        \PKGCnt[6]_net_1\, Y => \ByteDout_RNO_2[3]_net_1\);
    
    \CRC_Reg_RNO_2[5]\ : NOR2A
      port map(A => N_690_0, B => \CRC_Reg[4]_net_1\, Y => N_612);
    
    \Din_Delay4_RNIR778[1]\ : MX2
      port map(A => \Din_Delay4[1]_net_1\, B => 
        \CRC_Reg[33]_net_1\, S => \CRC_ResultAva\, Y => N_423);
    
    \CRC_Reg[28]\ : DFN1C0
      port map(D => N_23, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \CRC_Reg[28]_net_1\);
    
    \CRC_Reg_RNO[15]\ : NOR3
      port map(A => N_443, B => \CRC_Reg_14_2_i_0[15]\, C => 
        N_688, Y => N_290);
    
    \CRC_Reg_RNO_1[13]\ : OAI1
      port map(A => \CRC_Reg[5]_net_1\, B => N_692_0, C => 
        CMOS_DrvX_0_LVDSen_0, Y => \CRC_Reg_14_2_i_0[13]\);
    
    \PKGCnt[3]\ : DFN1E0C0
      port map(D => N_397_i_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => N_329_0, Q => 
        \PKGCnt[3]_net_1\);
    
    \DataClkCnt_RNI11SF[4]\ : NOR2B
      port map(A => N_305, B => \DataClkCnt[4]_net_1\, Y => N_309);
    
    \CRC_Reg_RNO_1[10]\ : OAI1
      port map(A => \CRC_Reg[2]_net_1\, B => N_692, C => 
        CMOS_DrvX_0_LVDSen_1, Y => \CRC_Reg_14_i_0_0[10]\);
    
    \CRC_Reg_RNO_1[1]\ : NOR2
      port map(A => N_450, B => \ByteDout[1]_net_1\, Y => N_623);
    
    \Prstate_RNO[2]\ : AO1C
      port map(A => \ClkEn_0\, B => \Prstate_ns_0_a5_0[5]\, C => 
        N_548, Y => \Prstate_ns[5]\);
    
    un1_clkdivcnt_I_13 : XOR2
      port map(A => N_4, B => \ClkDivCnt[3]_net_1\, Y => I_13);
    
    \DelayCnt_RNIL3IL[3]\ : AO1C
      port map(A => N_698, B => \DelayCnt[3]_net_1\, C => N_1049, 
        Y => N_335);
    
    \PKGCnt[15]\ : DFN1E0C0
      port map(D => PKGCnt_n15, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => N_329_0, Q => 
        \PKGCnt[15]_net_1\);
    
    \DataClkCnt_RNO[7]\ : NOR3A
      port map(A => N_979, B => N_990, C => N_992, Y => N_28);
    
    ClkEn_0_RNIF0SD : NOR2A
      port map(A => \ClkEn_0\, B => N_313, Y => N_333_i_0);
    
    \CRC_Reg[9]\ : DFN1C0
      port map(D => \CRC_Reg_RNO[9]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \CRC_Reg[9]_net_1\);
    
    \DataClkCnt_RNI4QG9[2]\ : NOR2B
      port map(A => N_298, B => \DataClkCnt[2]_net_1\, Y => N_302);
    
    \DataClkCnt[8]\ : DFN1C0
      port map(D => DataClkCnt_e8, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \DataClkCnt[8]_net_1\);
    
    \ByteDout_RNO_9[0]\ : NOR2B
      port map(A => \PKGCnt[3]_net_1\, B => DelayCnt_c0, Y => 
        \ByteDout_8_1_a5_3_0[0]\);
    
    \CRC_Reg_RNO_0[22]\ : AO1C
      port map(A => \CRC_Reg[21]_net_1\, B => N_690_0, C => 
        CMOS_DrvX_0_LVDSen_0, Y => \CRC_Reg_14_2_i_0[22]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \CRC_Reg[11]\ : DFN1C0
      port map(D => N_11, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \CRC_Reg[11]_net_1\);
    
    \Din_Delay4[2]\ : DFN1E1P0
      port map(D => \Din_Delay3[2]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, PRE => PLL_Test1_0_SysRst_O, E
         => \ClkEn\, Q => \Din_Delay4[2]_net_1\);
    
    \ByteDout_RNO_5[3]\ : OA1A
      port map(A => \Prstate[4]_net_1\, B => \Fifo_dout[3]\, C
         => N_1049, Y => \ByteDout_8_i_0[3]\);
    
    \ByteDout_RNO_3[4]\ : NOR3C
      port map(A => \ByteDout_RNO_4[4]_net_1\, B => 
        \ByteDout_RNO_5[4]_net_1\, C => N_1055, Y => 
        \ByteDout_8_i_1[4]\);
    
    \DelayCnt_RNI1M8L[2]\ : OR3A
      port map(A => \DelayCnt[2]_net_1\, B => N_313, C => N_693, 
        Y => N_705);
    
    CRC_ResultAva_RNO_1 : NOR2
      port map(A => \DelayCnt[1]_net_1\, B => \DelayCnt[3]_net_1\, 
        Y => CRC_ResultAva_3_0_a5_0_1);
    
    \StepCnt[3]\ : DFN1E1P0
      port map(D => N_211, CLK => PLL_Test1_0_Sys_66M_Clk, PRE
         => PLL_Test1_0_SysRst_O, E => StepCnte, Q => 
        \StepCnt[3]_net_1\);
    
    DataOk : DFN1E1C0
      port map(D => DataOk_0_sqmuxa, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => \ClkEn_1\, Q => \DataOk\);
    
    \ByteDout_RNO_4[6]\ : OA1A
      port map(A => \DelayCnt[3]_net_1\, B => N_698, C => 
        \ByteDout_RNO_8[6]_net_1\, Y => \ByteDout_8_i_2[6]\);
    
    \CRC_Reg_RNO[4]\ : OA1B
      port map(A => \CRC_Reg[4]_net_1\, B => N_448, C => 
        \CRC_Reg_14_i_0_1[4]\, Y => \CRC_Reg_RNO[4]_net_1\);
    
    \DataClkCnt_RNO[11]\ : AO1B
      port map(A => N_363, B => \DataClkCnt[11]_net_1\, C => 
        DataClkCnt_e11_0_0_0, Y => DataClkCnt_e11);
    
    \DataClkCnt_RNIMKIC[7]\ : NOR3C
      port map(A => \DataClkCnt[10]_net_1\, B => 
        \DataClkCnt[7]_net_1\, C => DataOk_0_sqmuxa_0_a2_0_a5_4, 
        Y => DataOk_0_sqmuxa_0_a2_0_a5_8);
    
    \ByteDout[7]\ : DFN1E1P0
      port map(D => N_186_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        PRE => PLL_Test1_0_SysRst_O, E => N_721, Q => 
        \ByteDout[7]_net_1\);
    
    \CRC_Reg_RNO[21]\ : OA1B
      port map(A => \CRC_Reg[21]_net_1\, B => N_291_0, C => 
        \CRC_Reg_14_2_i_1[21]\, Y => N_226);
    
    \ByteDout_RNO_0[0]\ : NOR3C
      port map(A => \ByteDout_8_1_2[0]\, B => \ByteDout_8_1_1[0]\, 
        C => N_1033, Y => \ByteDout_8_1_4[0]\);
    
    \ByteDout_RNO_2[6]\ : NOR3B
      port map(A => \ByteDout_8_i_1[6]\, B => \ByteDout_8_i_2[6]\, 
        C => N_708, Y => \ByteDout_8_i_4[6]\);
    
    \ByteDout_RNO_0[6]\ : OR2
      port map(A => \rowcnt[6]_net_1\, B => N_705, Y => 
        \ByteDout_RNO_0[6]_net_1\);
    
    \PKGCnt_RNO[3]\ : XNOR2
      port map(A => \PKGCnt[3]_net_1\, B => N_295, Y => 
        N_397_i_i_0);
    
    \CRC_Reg_RNO[20]\ : NOR3
      port map(A => N_432, B => \CRC_Reg_14_2_i_0[20]\, C => 
        N_597, Y => N_240);
    
    \ByteDout_RNO_6[7]\ : OR2A
      port map(A => \Prstate[4]_net_1\, B => \Fifo_dout[7]\, Y
         => \ByteDout_RNO_6[7]_net_1\);
    
    \ByteDout_RNO_3[0]\ : OR3B
      port map(A => N_412, B => \DelayCnt[1]_net_1\, C => N_698, 
        Y => N_1033);
    
    \ByteDout_RNO_2[4]\ : OA1
      port map(A => N_705, B => \rowcnt[4]_net_1\, C => 
        \ByteDout_8_i_1[4]\, Y => \ByteDout_8_i_3[4]\);
    
    \StepCnt[1]\ : DFN1E1C0
      port map(D => N_6, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => StepCnte, Q => 
        \StepCnt[1]_net_1\);
    
    \rowcnt_RNO[1]\ : XOR2
      port map(A => \rowcnt[1]_net_1\, B => \rowcnt[0]_net_1\, Y
         => N_385_i);
    
    \FrameCnt[8]\ : DFN1E0C0
      port map(D => N_446_i_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => N_365, Q => 
        \FrameCnt[8]_net_1\);
    
    \FrameCnt[6]\ : DFN1E0C0
      port map(D => N_415_i_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => N_365, Q => 
        \FrameCnt[6]_net_1\);
    
    \CRC_Reg_RNO_0[6]\ : AO1D
      port map(A => N_450, B => \ByteDout[6]_net_1\, C => N_609, 
        Y => \CRC_Reg_14_i_0_0[6]\);
    
    ClkEn_1_RNIHLPK : OR2A
      port map(A => N_450, B => N_690, Y => N_448);
    
    \CRC_Reg_RNO_0[39]\ : AO1D
      port map(A => N_692_0, B => \CRC_Reg[31]_net_1\, C => 
        \CRC_Reg_14_2_i_0[39]\, Y => \CRC_Reg_14_2_i_1[39]\);
    
    \Shifter_RNO[4]\ : MX2
      port map(A => \Shifter[5]_net_1\, B => \TenbitDout[4]\, S
         => \PtS_En\, Y => \Shifter_4[4]\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3;
use proasic3.all;

entity My_adder0_1 is

    port( intData2acc_RNIEVV9                         : in    std_logic_vector(64 to 64);
          intData2acc_RNIDVV9                         : in    std_logic_vector(63 to 63);
          intData2acc_RNIGVV9                         : in    std_logic_vector(66 to 66);
          intData2acc_RNIDRV9                         : in    std_logic_vector(56 to 56);
          intData2acc_RNIERV9                         : in    std_logic_vector(57 to 57);
          intData2acc_RNIHVV9                         : in    std_logic_vector(67 to 67);
          intData2acc_RNIAVV9                         : in    std_logic_vector(60 to 60);
          intData2acc_RNIBVV9                         : in    std_logic_vector(61 to 61);
          intData2acc_RNIFVV9                         : in    std_logic_vector(65 to 65);
          intData2acc_RNIPB46                         : in    std_logic_vector(71 to 71);
          intData2acc_RNIGRV9                         : in    std_logic_vector(59 downto 58);
          intData2acc_RNICVV9                         : in    std_logic_vector(62 to 62);
          intData2acc_RNID30A                         : in    std_logic_vector(70 to 70);
          intData2acc_RNIARV9                         : in    std_logic_vector(54 to 54);
          intData2acc_RNIBRV9                         : in    std_logic_vector(55 to 55);
          \Z\\My_adder0_3_Sum_[15]\\\                 : out   std_logic;
          \Z\\My_adder0_3_Sum_[12]\\\                 : out   std_logic;
          \Z\\My_adder0_3_Sum_[6]\\\                  : out   std_logic;
          \Z\\My_adder0_3_Sum_[10]\\\                 : out   std_logic;
          \Z\\My_adder0_3_Sum_[9]\\\                  : out   std_logic;
          \Z\\My_adder0_3_Sum_[7]\\\                  : out   std_logic;
          N_6                                         : in    std_logic;
          \Z\\My_adder0_3_Sum_[11]\\\                 : out   std_logic;
          \Z\\My_adder0_3_Sum_[1]\\\                  : out   std_logic;
          \Z\\My_adder0_3_Sum_[3]\\\                  : out   std_logic;
          \Z\\My_adder0_3_Sum_[13]\\\                 : out   std_logic;
          \Z\\My_adder0_3_Sum_[0]\\\                  : out   std_logic;
          \Z\\My_adder0_3_Sum_[8]\\\                  : out   std_logic;
          \Z\\My_adder0_3_Sum_[14]\\\                 : out   std_logic;
          \Z\\My_adder0_3_Sum_[2]\\\                  : out   std_logic;
          \Z\\My_adder0_3_Sum_[4]\\\                  : out   std_logic;
          N_4                                         : in    std_logic;
          \Z\\My_adder0_3_Sum_[5]\\\                  : out   std_logic;
          \Z\\My_adder0_3_Sum_[17]\\\                 : out   std_logic;
          My_adder0_1_GND                             : in    std_logic;
          \Z\\My_adder0_3_Sum_[16]\\\                 : out   std_logic;
          \Z\\adc_muxtmp_test_0_DataOut55to42_[43]\\\ : in    std_logic
        );

end My_adder0_1;

architecture DEF_ARCH of My_adder0_1 is 

  component XOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MAJ3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component AND2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal Carry_1_net, Carry_0_net, Carry_15_net, Carry_8_net, 
        Carry_7_net, Carry_5_net, Carry_4_net, Carry_16_net, 
        Carry_11_net, Carry_10_net, Carry_6_net, Carry_13_net, 
        Carry_12_net, Carry_3_net, Carry_2_net, Carry_14_net, 
        Carry_9_net, \GND\, \VCC\, GND_0, VCC_0 : std_logic;

begin 


    XOR3_Sum_16_inst : XOR3
      port map(A => My_adder0_1_GND, B => intData2acc_RNID30A(70), 
        C => Carry_15_net, Y => \Z\\My_adder0_3_Sum_[16]\\\);
    
    MAJ3_Carry_8_inst : MAJ3
      port map(A => Carry_7_net, B => My_adder0_1_GND, C => 
        intData2acc_RNICVV9(62), Y => Carry_8_net);
    
    MAJ3_Carry_9_inst : MAJ3
      port map(A => Carry_8_net, B => My_adder0_1_GND, C => 
        intData2acc_RNIDVV9(63), Y => Carry_9_net);
    
    XOR3_Sum_5_inst : XOR3
      port map(A => My_adder0_1_GND, B => intData2acc_RNIGRV9(59), 
        C => Carry_4_net, Y => \Z\\My_adder0_3_Sum_[5]\\\);
    
    XOR3_Sum_2_inst : XOR3
      port map(A => My_adder0_1_GND, B => intData2acc_RNIDRV9(56), 
        C => Carry_1_net, Y => \Z\\My_adder0_3_Sum_[2]\\\);
    
    XOR3_Sum_4_inst : XOR3
      port map(A => My_adder0_1_GND, B => intData2acc_RNIGRV9(58), 
        C => Carry_3_net, Y => \Z\\My_adder0_3_Sum_[4]\\\);
    
    XOR3_Sum_11_inst : XOR3
      port map(A => My_adder0_1_GND, B => intData2acc_RNIFVV9(65), 
        C => Carry_10_net, Y => \Z\\My_adder0_3_Sum_[11]\\\);
    
    XOR3_Sum_12_inst : XOR3
      port map(A => My_adder0_1_GND, B => intData2acc_RNIGVV9(66), 
        C => Carry_11_net, Y => \Z\\My_adder0_3_Sum_[12]\\\);
    
    MAJ3_Carry_5_inst : MAJ3
      port map(A => Carry_4_net, B => My_adder0_1_GND, C => 
        intData2acc_RNIGRV9(59), Y => Carry_5_net);
    
    MAJ3_Carry_2_inst : MAJ3
      port map(A => Carry_1_net, B => My_adder0_1_GND, C => 
        intData2acc_RNIDRV9(56), Y => Carry_2_net);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    MAJ3_Carry_4_inst : MAJ3
      port map(A => Carry_3_net, B => My_adder0_1_GND, C => 
        intData2acc_RNIGRV9(58), Y => Carry_4_net);
    
    XOR3_Sum_13_inst : XOR3
      port map(A => My_adder0_1_GND, B => intData2acc_RNIHVV9(67), 
        C => Carry_12_net, Y => \Z\\My_adder0_3_Sum_[13]\\\);
    
    AND2_Carry_0_inst_RNI9VHF : MAJ3
      port map(A => Carry_0_net, B => 
        \Z\\adc_muxtmp_test_0_DataOut55to42_[43]\\\, C => 
        intData2acc_RNIBRV9(55), Y => Carry_1_net);
    
    XOR3_Sum_1_inst : XOR3
      port map(A => \Z\\adc_muxtmp_test_0_DataOut55to42_[43]\\\, 
        B => intData2acc_RNIBRV9(55), C => Carry_0_net, Y => 
        \Z\\My_adder0_3_Sum_[1]\\\);
    
    MAJ3_Carry_12_inst : MAJ3
      port map(A => Carry_11_net, B => My_adder0_1_GND, C => 
        intData2acc_RNIGVV9(66), Y => Carry_12_net);
    
    XOR3_Sum_17_inst : XOR3
      port map(A => My_adder0_1_GND, B => intData2acc_RNIPB46(71), 
        C => Carry_16_net, Y => \Z\\My_adder0_3_Sum_[17]\\\);
    
    MAJ3_Carry_7_inst : MAJ3
      port map(A => Carry_6_net, B => My_adder0_1_GND, C => 
        intData2acc_RNIBVV9(61), Y => Carry_7_net);
    
    GND_i : GND
      port map(Y => \GND\);
    
    XOR3_Sum_6_inst : XOR3
      port map(A => My_adder0_1_GND, B => intData2acc_RNIAVV9(60), 
        C => Carry_5_net, Y => \Z\\My_adder0_3_Sum_[6]\\\);
    
    MAJ3_Carry_14_inst : MAJ3
      port map(A => Carry_13_net, B => My_adder0_1_GND, C => N_4, 
        Y => Carry_14_net);
    
    MAJ3_Carry_13_inst : MAJ3
      port map(A => Carry_12_net, B => My_adder0_1_GND, C => 
        intData2acc_RNIHVV9(67), Y => Carry_13_net);
    
    XOR3_Sum_3_inst : XOR3
      port map(A => My_adder0_1_GND, B => intData2acc_RNIERV9(57), 
        C => Carry_2_net, Y => \Z\\My_adder0_3_Sum_[3]\\\);
    
    XOR3_Sum_14_inst : XOR3
      port map(A => My_adder0_1_GND, B => N_4, C => Carry_13_net, 
        Y => \Z\\My_adder0_3_Sum_[14]\\\);
    
    XOR3_Sum_8_inst : XOR3
      port map(A => My_adder0_1_GND, B => intData2acc_RNICVV9(62), 
        C => Carry_7_net, Y => \Z\\My_adder0_3_Sum_[8]\\\);
    
    MAJ3_Carry_11_inst : MAJ3
      port map(A => Carry_10_net, B => My_adder0_1_GND, C => 
        intData2acc_RNIFVV9(65), Y => Carry_11_net);
    
    MAJ3_Carry_16_inst : MAJ3
      port map(A => Carry_15_net, B => My_adder0_1_GND, C => 
        intData2acc_RNID30A(70), Y => Carry_16_net);
    
    XOR3_Sum_7_inst : XOR3
      port map(A => My_adder0_1_GND, B => intData2acc_RNIBVV9(61), 
        C => Carry_6_net, Y => \Z\\My_adder0_3_Sum_[7]\\\);
    
    MAJ3_Carry_10_inst : MAJ3
      port map(A => Carry_9_net, B => My_adder0_1_GND, C => 
        intData2acc_RNIEVV9(64), Y => Carry_10_net);
    
    MAJ3_Carry_3_inst : MAJ3
      port map(A => Carry_2_net, B => My_adder0_1_GND, C => 
        intData2acc_RNIERV9(57), Y => Carry_3_net);
    
    XOR3_Sum_15_inst : XOR3
      port map(A => My_adder0_1_GND, B => N_6, C => Carry_14_net, 
        Y => \Z\\My_adder0_3_Sum_[15]\\\);
    
    AND2_Carry_0_inst : AND2
      port map(A => \Z\\adc_muxtmp_test_0_DataOut55to42_[43]\\\, 
        B => intData2acc_RNIARV9(54), Y => Carry_0_net);
    
    MAJ3_Carry_15_inst : MAJ3
      port map(A => Carry_14_net, B => My_adder0_1_GND, C => N_6, 
        Y => Carry_15_net);
    
    XOR3_Sum_9_inst : XOR3
      port map(A => My_adder0_1_GND, B => intData2acc_RNIDVV9(63), 
        C => Carry_8_net, Y => \Z\\My_adder0_3_Sum_[9]\\\);
    
    XOR2_Sum_0_inst : XOR2
      port map(A => \Z\\adc_muxtmp_test_0_DataOut55to42_[43]\\\, 
        B => intData2acc_RNIARV9(54), Y => 
        \Z\\My_adder0_3_Sum_[0]\\\);
    
    MAJ3_Carry_6_inst : MAJ3
      port map(A => Carry_5_net, B => My_adder0_1_GND, C => 
        intData2acc_RNIAVV9(60), Y => Carry_6_net);
    
    XOR3_Sum_10_inst : XOR3
      port map(A => My_adder0_1_GND, B => intData2acc_RNIEVV9(64), 
        C => Carry_9_net, Y => \Z\\My_adder0_3_Sum_[10]\\\);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3;
use proasic3.all;

entity Fifo_rd is

    port( \Z\\Fifo_wr_0_Q_[27]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[23]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[69]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[1]\\\              : out   std_logic;
          \Z\\Fifo_wr_0_Q_[67]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[4]\\\              : out   std_logic;
          \Z\\Fifo_wr_0_Q_[63]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[7]\\\              : out   std_logic;
          \Z\\Fifo_wr_0_Q_[56]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[25]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[24]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[48]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[65]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[64]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[51]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[38]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[71]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[50]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[70]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[18]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[6]\\\              : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[71]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[70]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[69]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[68]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[67]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[66]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[65]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[64]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[63]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[62]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[61]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[60]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[59]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[58]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[57]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[56]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[55]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[54]\\\ : in    std_logic;
          \Z\\Fifo_wr_0_Q_[46]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[52]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[36]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[59]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[0]\\\              : out   std_logic;
          \Z\\Fifo_wr_0_Q_[16]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[57]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[41]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[53]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[40]\\\             : out   std_logic;
          Sdram_cmd_0_WFifo_re                : in    std_logic;
          \Z\\Fifo_wr_0_Q_[31]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[28]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[30]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[42]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[11]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[10]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[55]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[68]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[54]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[49]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[9]\\\              : out   std_logic;
          \Z\\Fifo_wr_0_Q_[5]\\\              : out   std_logic;
          Fifo_wr_0_AFULL                     : out   std_logic;
          \Z\\Fifo_wr_0_Q_[32]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[47]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[43]\\\             : out   std_logic;
          Main_ctl4SD_0_fifo_rst_n_3          : in    std_logic;
          \Z\\Fifo_wr_0_Q_[12]\\\             : out   std_logic;
          Main_ctl4SD_0_Fifo_wr               : in    std_logic;
          \Z\\Fifo_wr_0_Q_[26]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[39]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[19]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[37]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[3]\\\              : out   std_logic;
          \Z\\Fifo_wr_0_Q_[33]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[66]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[17]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[13]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[45]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[44]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[21]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[2]\\\              : out   std_logic;
          \Z\\Fifo_wr_0_Q_[20]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[61]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[35]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[34]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[60]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[15]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[14]\\\             : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[35]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[34]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[33]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[32]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[31]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[30]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[29]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[28]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[27]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[26]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[25]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[24]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[23]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[22]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[21]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[20]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[19]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[18]\\\ : in    std_logic;
          Main_ctl4SD_0_fifo_rst_n_4          : in    std_logic;
          \Z\\Fifo_wr_0_Q_[22]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[8]\\\              : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[53]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[52]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[51]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[50]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[49]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[48]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[47]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[46]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[45]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[44]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[43]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[42]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[41]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[40]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[39]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[38]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[37]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[36]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[17]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[16]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[15]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[14]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[13]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[12]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[11]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[10]\\\ : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[9]\\\  : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[8]\\\  : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[7]\\\  : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[6]\\\  : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[5]\\\  : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[4]\\\  : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[3]\\\  : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[2]\\\  : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[1]\\\  : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[0]\\\  : in    std_logic;
          Fifo_rd_VCC                         : in    std_logic;
          Main_ctl4SD_0_fifo_rst_n            : in    std_logic;
          \Z\\Fifo_wr_0_Q_[62]\\\             : out   std_logic;
          Main_ctl4SD_0_fifo_rst_n_5          : in    std_logic;
          \Z\\Fifo_wr_0_Q_[29]\\\             : out   std_logic;
          Main_ctl4SD_0_fifo_rst_n_6          : in    std_logic;
          PLL_Test1_0_Sys_66M_Clk             : in    std_logic;
          \Z\\Fifo_wr_0_Q_[58]\\\             : out   std_logic;
          Fifo_rd_GND                         : in    std_logic
        );

end Fifo_rd;

architecture DEF_ARCH of Fifo_rd is 

  component INV
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XNOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component BUFF
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component RAM512X18
    generic (MEMORYFILE:string := "");

    port( RADDR8 : in    std_logic := 'U';
          RADDR7 : in    std_logic := 'U';
          RADDR6 : in    std_logic := 'U';
          RADDR5 : in    std_logic := 'U';
          RADDR4 : in    std_logic := 'U';
          RADDR3 : in    std_logic := 'U';
          RADDR2 : in    std_logic := 'U';
          RADDR1 : in    std_logic := 'U';
          RADDR0 : in    std_logic := 'U';
          WADDR8 : in    std_logic := 'U';
          WADDR7 : in    std_logic := 'U';
          WADDR6 : in    std_logic := 'U';
          WADDR5 : in    std_logic := 'U';
          WADDR4 : in    std_logic := 'U';
          WADDR3 : in    std_logic := 'U';
          WADDR2 : in    std_logic := 'U';
          WADDR1 : in    std_logic := 'U';
          WADDR0 : in    std_logic := 'U';
          WD17   : in    std_logic := 'U';
          WD16   : in    std_logic := 'U';
          WD15   : in    std_logic := 'U';
          WD14   : in    std_logic := 'U';
          WD13   : in    std_logic := 'U';
          WD12   : in    std_logic := 'U';
          WD11   : in    std_logic := 'U';
          WD10   : in    std_logic := 'U';
          WD9    : in    std_logic := 'U';
          WD8    : in    std_logic := 'U';
          WD7    : in    std_logic := 'U';
          WD6    : in    std_logic := 'U';
          WD5    : in    std_logic := 'U';
          WD4    : in    std_logic := 'U';
          WD3    : in    std_logic := 'U';
          WD2    : in    std_logic := 'U';
          WD1    : in    std_logic := 'U';
          WD0    : in    std_logic := 'U';
          RW0    : in    std_logic := 'U';
          RW1    : in    std_logic := 'U';
          WW0    : in    std_logic := 'U';
          WW1    : in    std_logic := 'U';
          PIPE   : in    std_logic := 'U';
          REN    : in    std_logic := 'U';
          WEN    : in    std_logic := 'U';
          RCLK   : in    std_logic := 'U';
          WCLK   : in    std_logic := 'U';
          RESET  : in    std_logic := 'U';
          RD17   : out   std_logic;
          RD16   : out   std_logic;
          RD15   : out   std_logic;
          RD14   : out   std_logic;
          RD13   : out   std_logic;
          RD12   : out   std_logic;
          RD11   : out   std_logic;
          RD10   : out   std_logic;
          RD9    : out   std_logic;
          RD8    : out   std_logic;
          RD7    : out   std_logic;
          RD6    : out   std_logic;
          RD5    : out   std_logic;
          RD4    : out   std_logic;
          RD3    : out   std_logic;
          RD2    : out   std_logic;
          RD1    : out   std_logic;
          RD0    : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component NAND3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NAND2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal DVLDI_2, DVLDI, DVLDI_1, DVLDI_0, AND2_25_Y, AND3_1_Y, 
        XNOR2_6_Y, AND2_28_Y, MEM_RADDR_0_net, MEMORYRE, 
        XNOR2_8_Y, MEM_RADDR_3_net, WBINNXTSHIFT_3_net, XOR2_36_Y, 
        MEM_RADDR_4_net, QXI_58_net, QXI_29_net, 
        RBINNXTSHIFT_2_net, XOR2_10_Y, AO1_8_Y, QXI_62_net, 
        QXI_0_net, QXI_1_net, QXI_2_net, QXI_3_net, QXI_4_net, 
        QXI_5_net, QXI_6_net, QXI_7_net, QXI_8_net, QXI_9_net, 
        QXI_10_net, QXI_11_net, QXI_12_net, QXI_13_net, 
        QXI_14_net, QXI_15_net, QXI_16_net, QXI_17_net, 
        MEM_RADDR_1_net, MEM_RADDR_2_net, MEMRENEG, 
        MEM_WADDR_0_net, MEM_WADDR_1_net, MEM_WADDR_2_net, 
        MEM_WADDR_3_net, MEMWENEG, AO1_4_Y, XOR2_11_Y, AO1_0_Y, 
        AND2_3_Y, NAND2_1_Y, DFN1P0_EMPTY_1, XOR2_0_Y, 
        WBINNXTSHIFT_1_net, AND2_8_Y, AND2_21_Y, QXI_36_net, 
        QXI_37_net, QXI_38_net, QXI_39_net, QXI_40_net, 
        QXI_41_net, QXI_42_net, QXI_43_net, QXI_44_net, 
        QXI_45_net, QXI_46_net, QXI_47_net, QXI_48_net, 
        QXI_49_net, QXI_50_net, QXI_51_net, QXI_52_net, 
        QXI_53_net, QXI_22_net, RBINNXTSHIFT_0_net, QXI_18_net, 
        QXI_19_net, QXI_20_net, QXI_21_net, QXI_23_net, 
        QXI_24_net, QXI_25_net, QXI_26_net, QXI_27_net, 
        QXI_28_net, QXI_30_net, QXI_31_net, QXI_32_net, 
        QXI_33_net, QXI_34_net, QXI_35_net, XOR2_28_Y, QXI_60_net, 
        RBINNXTSHIFT_1_net, XOR2_29_Y, QXI_61_net, XOR2_3_Y, 
        INV_2_Y, MEMORYWE, WDIFF_4_net, XOR2_21_Y, AO1_6_Y, 
        AO1_5_Y, AND2_24_Y, AO1_11_Y, XNOR2_5_Y, FULLINT, 
        AND2_7_Y, XOR2_23_Y, AND2_4_Y, XNOR2_7_Y, OR2A_0_Y, 
        WDIFF_2_net, AO1_13_Y, XOR2_4_Y, NOR2A_0_Y, 
        WBINNXTSHIFT_0_net, AND2_17_Y, INV_3_Y, QXI_66_net, 
        EMPTYINT, XOR2_35_Y, AO1_10_Y, AND2_1_Y, AOI1_0_Y, 
        AND2_6_Y, NAND3A_1_Y, NOR3_0_Y, OA1A_0_Y, WDIFF_3_net, 
        WDIFF_1_net, XOR2_14_Y, AND2A_0_Y, XOR2_2_Y, XOR2_18_Y, 
        AND2_18_Y, NAND2_0_Y, XNOR2_10_Y, RBINNXTSHIFT_4_net, 
        MEM_WADDR_4_net, AND2A_1_Y, DFN1C0_FULL_1, NOR3A_0_Y, 
        NAND3A_0_Y, OR2_0_Y, OR2A_1_Y, AO1C_0_Y, WDIFF_0_net, 
        AND2_9_Y, QXI_54_net, OR3_0_Y, AND2_22_Y, AND2_2_Y, 
        QXI_68_net, QXI_55_net, XOR2_32_Y, RBINNXTSHIFT_3_net, 
        AO1_7_Y, XNOR2_3_Y, INV_1_Y, XOR2_7_Y, WBINNXTSHIFT_2_net, 
        INV_4_Y, XNOR2_1_Y, AND2_13_Y, XOR2_9_Y, AO1_3_Y, 
        AND2_12_Y, QXI_57_net, XOR2_13_Y, QXI_59_net, XNOR2_4_Y, 
        XOR2_20_Y, OA1C_0_Y, WBINNXTSHIFT_4_net, XOR2_16_Y, 
        QXI_56_net, QXI_63_net, QXI_64_net, QXI_65_net, 
        QXI_67_net, QXI_69_net, QXI_70_net, QXI_71_net, AND2_31_Y, 
        XNOR2_0_Y, XOR2_1_Y, XNOR2_2_Y, AND3_0_Y, XNOR2_9_Y, 
        INV_0_Y, \GND\, \VCC\, GND_0, VCC_0 : std_logic;

begin 


    INV_0 : INV
      port map(A => MEM_RADDR_4_net, Y => INV_0_Y);
    
    NOR3_0 : NOR3
      port map(A => OA1A_0_Y, B => AND2A_0_Y, C => OA1C_0_Y, Y
         => NOR3_0_Y);
    
    AND2_2 : AND2
      port map(A => INV_1_Y, B => INV_3_Y, Y => AND2_2_Y);
    
    DFN1E1C0_Q_27_inst : DFN1E1C0
      port map(D => QXI_27_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_5, E => DVLDI_0, Q => 
        \Z\\Fifo_wr_0_Q_[27]\\\);
    
    AO1_11 : AO1
      port map(A => XOR2_1_Y, B => AND2_4_Y, C => AND2_21_Y, Y
         => AO1_11_Y);
    
    AND2_22 : AND2
      port map(A => WBINNXTSHIFT_1_net, B => INV_1_Y, Y => 
        AND2_22_Y);
    
    XNOR2_9 : XNOR2
      port map(A => MEM_RADDR_2_net, B => WBINNXTSHIFT_2_net, Y
         => XNOR2_9_Y);
    
    DFN1C0_FULL : DFN1C0
      port map(D => FULLINT, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => Main_ctl4SD_0_fifo_rst_n_4, Q => DFN1C0_FULL_1);
    
    DFN1E1C0_Q_37_inst : DFN1E1C0
      port map(D => QXI_37_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_5, E => DVLDI_1, Q => 
        \Z\\Fifo_wr_0_Q_[37]\\\);
    
    DFN1E1C0_Q_23_inst : DFN1E1C0
      port map(D => QXI_23_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_5, E => DVLDI_0, Q => 
        \Z\\Fifo_wr_0_Q_[23]\\\);
    
    XOR2_23 : XOR2
      port map(A => MEM_RADDR_4_net, B => WBINNXTSHIFT_4_net, Y
         => XOR2_23_Y);
    
    XOR2_1 : XOR2
      port map(A => MEM_RADDR_3_net, B => Fifo_rd_GND, Y => 
        XOR2_1_Y);
    
    DFN1E1C0_Q_54_inst : DFN1E1C0
      port map(D => QXI_54_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_6, E => DVLDI_2, Q => 
        \Z\\Fifo_wr_0_Q_[54]\\\);
    
    DFN1E1C0_Q_33_inst : DFN1E1C0
      port map(D => QXI_33_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_5, E => DVLDI_1, Q => 
        \Z\\Fifo_wr_0_Q_[33]\\\);
    
    INV_1 : INV
      port map(A => MEM_RADDR_1_net, Y => INV_1_Y);
    
    AO1_7 : AO1
      port map(A => XOR2_7_Y, B => OR3_0_Y, C => AND2_31_Y, Y => 
        AO1_7_Y);
    
    AND2_18 : AND2
      port map(A => MEM_WADDR_1_net, B => Fifo_rd_GND, Y => 
        AND2_18_Y);
    
    DFN1C0_MEM_WADDR_2_inst : DFN1C0
      port map(D => WBINNXTSHIFT_2_net, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => 
        Main_ctl4SD_0_fifo_rst_n_4, Q => MEM_WADDR_2_net);
    
    AND2_1 : AND2
      port map(A => MEM_WADDR_3_net, B => Fifo_rd_GND, Y => 
        AND2_1_Y);
    
    AO1_8 : AO1
      port map(A => XOR2_2_Y, B => AND2_28_Y, C => AND2_13_Y, Y
         => AO1_8_Y);
    
    DFN1E1C0_Q_61_inst : DFN1E1C0
      port map(D => QXI_61_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_6, E => DVLDI_2, Q => 
        \Z\\Fifo_wr_0_Q_[61]\\\);
    
    XOR2_20 : XOR2
      port map(A => WBINNXTSHIFT_2_net, B => INV_4_Y, Y => 
        XOR2_20_Y);
    
    DFN1E1C0_Q_2_inst : DFN1E1C0
      port map(D => QXI_2_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_5, E => DVLDI_0, Q => 
        \Z\\Fifo_wr_0_Q_[2]\\\);
    
    AND2_7 : AND2
      port map(A => AND3_0_Y, B => XNOR2_8_Y, Y => AND2_7_Y);
    
    DFN1C0_DVLDI_RNI1QG2_0 : BUFF
      port map(A => DVLDI, Y => DVLDI_0);
    
    AND2_12 : AND2
      port map(A => XOR2_11_Y, B => XOR2_35_Y, Y => AND2_12_Y);
    
    AND2A_1 : AND2A
      port map(A => DFN1P0_EMPTY_1, B => Sdram_cmd_0_WFifo_re, Y
         => AND2A_1_Y);
    
    DFN1E1C0_Q_65_inst : DFN1E1C0
      port map(D => QXI_65_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n, E => DVLDI_2, Q => 
        \Z\\Fifo_wr_0_Q_[65]\\\);
    
    AND2_EMPTYINT : AND2
      port map(A => AND2_25_Y, B => XNOR2_10_Y, Y => EMPTYINT);
    
    RAM512X18_QXI_17_inst : RAM512X18
      port map(RADDR8 => Fifo_rd_GND, RADDR7 => Fifo_rd_GND, 
        RADDR6 => Fifo_rd_GND, RADDR5 => Fifo_rd_GND, RADDR4 => 
        Fifo_rd_GND, RADDR3 => MEM_RADDR_3_net, RADDR2 => 
        MEM_RADDR_2_net, RADDR1 => MEM_RADDR_1_net, RADDR0 => 
        MEM_RADDR_0_net, WADDR8 => Fifo_rd_GND, WADDR7 => 
        Fifo_rd_GND, WADDR6 => Fifo_rd_GND, WADDR5 => Fifo_rd_GND, 
        WADDR4 => Fifo_rd_GND, WADDR3 => MEM_WADDR_3_net, WADDR2
         => MEM_WADDR_2_net, WADDR1 => MEM_WADDR_1_net, WADDR0
         => MEM_WADDR_0_net, WD17 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[17]\\\, WD16 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[16]\\\, WD15 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[15]\\\, WD14 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[14]\\\, WD13 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[13]\\\, WD12 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[12]\\\, WD11 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[11]\\\, WD10 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[10]\\\, WD9 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[9]\\\, WD8 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[8]\\\, WD7 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[7]\\\, WD6 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[6]\\\, WD5 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[5]\\\, WD4 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[4]\\\, WD3 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[3]\\\, WD2 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[2]\\\, WD1 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[1]\\\, WD0 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[0]\\\, RW0 => Fifo_rd_GND, 
        RW1 => Fifo_rd_VCC, WW0 => Fifo_rd_GND, WW1 => 
        Fifo_rd_VCC, PIPE => Fifo_rd_GND, REN => MEMRENEG, WEN
         => MEMWENEG, RCLK => PLL_Test1_0_Sys_66M_Clk, WCLK => 
        PLL_Test1_0_Sys_66M_Clk, RESET => 
        Main_ctl4SD_0_fifo_rst_n, RD17 => QXI_17_net, RD16 => 
        QXI_16_net, RD15 => QXI_15_net, RD14 => QXI_14_net, RD13
         => QXI_13_net, RD12 => QXI_12_net, RD11 => QXI_11_net, 
        RD10 => QXI_10_net, RD9 => QXI_9_net, RD8 => QXI_8_net, 
        RD7 => QXI_7_net, RD6 => QXI_6_net, RD5 => QXI_5_net, RD4
         => QXI_4_net, RD3 => QXI_3_net, RD2 => QXI_2_net, RD1
         => QXI_1_net, RD0 => QXI_0_net);
    
    DFN1C0_DVLDI_RNI1QG2_1 : BUFF
      port map(A => DVLDI, Y => DVLDI_2);
    
    XOR2_21 : XOR2
      port map(A => WBINNXTSHIFT_4_net, B => INV_0_Y, Y => 
        XOR2_21_Y);
    
    DFN1C0_MEM_RADDR_0_inst : DFN1C0
      port map(D => RBINNXTSHIFT_0_net, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => 
        Main_ctl4SD_0_fifo_rst_n_4, Q => MEM_RADDR_0_net);
    
    DFN1E1C0_Q_5_inst : DFN1E1C0
      port map(D => QXI_5_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_6, E => DVLDI_2, Q => 
        \Z\\Fifo_wr_0_Q_[5]\\\);
    
    DFN1E1C0_Q_14_inst : DFN1E1C0
      port map(D => QXI_14_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_4, E => DVLDI_0, Q => 
        \Z\\Fifo_wr_0_Q_[14]\\\);
    
    XOR2_16 : XOR2
      port map(A => MEM_WADDR_4_net, B => Fifo_rd_GND, Y => 
        XOR2_16_Y);
    
    DFN1E1C0_Q_66_inst : DFN1E1C0
      port map(D => QXI_66_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n, E => DVLDI_2, Q => 
        \Z\\Fifo_wr_0_Q_[66]\\\);
    
    RAM512X18_QXI_53_inst : RAM512X18
      port map(RADDR8 => Fifo_rd_GND, RADDR7 => Fifo_rd_GND, 
        RADDR6 => Fifo_rd_GND, RADDR5 => Fifo_rd_GND, RADDR4 => 
        Fifo_rd_GND, RADDR3 => MEM_RADDR_3_net, RADDR2 => 
        MEM_RADDR_2_net, RADDR1 => MEM_RADDR_1_net, RADDR0 => 
        MEM_RADDR_0_net, WADDR8 => Fifo_rd_GND, WADDR7 => 
        Fifo_rd_GND, WADDR6 => Fifo_rd_GND, WADDR5 => Fifo_rd_GND, 
        WADDR4 => Fifo_rd_GND, WADDR3 => MEM_WADDR_3_net, WADDR2
         => MEM_WADDR_2_net, WADDR1 => MEM_WADDR_1_net, WADDR0
         => MEM_WADDR_0_net, WD17 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[53]\\\, WD16 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[52]\\\, WD15 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[51]\\\, WD14 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[50]\\\, WD13 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[49]\\\, WD12 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[48]\\\, WD11 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[47]\\\, WD10 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[46]\\\, WD9 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[45]\\\, WD8 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[44]\\\, WD7 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[43]\\\, WD6 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[42]\\\, WD5 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[41]\\\, WD4 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[40]\\\, WD3 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[39]\\\, WD2 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[38]\\\, WD1 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[37]\\\, WD0 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[36]\\\, RW0 => Fifo_rd_GND, 
        RW1 => Fifo_rd_VCC, WW0 => Fifo_rd_GND, WW1 => 
        Fifo_rd_VCC, PIPE => Fifo_rd_GND, REN => MEMRENEG, WEN
         => MEMWENEG, RCLK => PLL_Test1_0_Sys_66M_Clk, WCLK => 
        PLL_Test1_0_Sys_66M_Clk, RESET => 
        Main_ctl4SD_0_fifo_rst_n, RD17 => QXI_53_net, RD16 => 
        QXI_52_net, RD15 => QXI_51_net, RD14 => QXI_50_net, RD13
         => QXI_49_net, RD12 => QXI_48_net, RD11 => QXI_47_net, 
        RD10 => QXI_46_net, RD9 => QXI_45_net, RD8 => QXI_44_net, 
        RD7 => QXI_43_net, RD6 => QXI_42_net, RD5 => QXI_41_net, 
        RD4 => QXI_40_net, RD3 => QXI_39_net, RD2 => QXI_38_net, 
        RD1 => QXI_37_net, RD0 => QXI_36_net);
    
    DFN1E1C0_Q_62_inst : DFN1E1C0
      port map(D => QXI_62_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n, E => DVLDI_2, Q => 
        \Z\\Fifo_wr_0_Q_[62]\\\);
    
    OR2_0 : OR2
      port map(A => AOI1_0_Y, B => DFN1C0_FULL_1, Y => OR2_0_Y);
    
    MEMWEBUBBLE : INV
      port map(A => MEMORYWE, Y => MEMWENEG);
    
    AND2_6 : AND2
      port map(A => XNOR2_4_Y, B => XNOR2_1_Y, Y => AND2_6_Y);
    
    AND3_0 : AND3
      port map(A => XNOR2_0_Y, B => XNOR2_7_Y, C => XNOR2_9_Y, Y
         => AND3_0_Y);
    
    DFN1E1C0_Q_0_inst : DFN1E1C0
      port map(D => QXI_0_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_4, E => DVLDI_0, Q => 
        \Z\\Fifo_wr_0_Q_[0]\\\);
    
    INV_3 : INV
      port map(A => NOR2A_0_Y, Y => INV_3_Y);
    
    XNOR2_2 : XNOR2
      port map(A => RBINNXTSHIFT_1_net, B => MEM_WADDR_1_net, Y
         => XNOR2_2_Y);
    
    DFN1E1C0_Q_29_inst : DFN1E1C0
      port map(D => QXI_29_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_5, E => DVLDI_0, Q => 
        \Z\\Fifo_wr_0_Q_[29]\\\);
    
    XOR2_WBINNXTSHIFT_2_inst : XOR2
      port map(A => XOR2_13_Y, B => AO1_0_Y, Y => 
        WBINNXTSHIFT_2_net);
    
    XOR2_4 : XOR2
      port map(A => MEM_RADDR_2_net, B => Fifo_rd_GND, Y => 
        XOR2_4_Y);
    
    AND3_1 : AND3
      port map(A => XNOR2_3_Y, B => XNOR2_2_Y, C => XNOR2_5_Y, Y
         => AND3_1_Y);
    
    AND2_24 : AND2
      port map(A => XOR2_4_Y, B => XOR2_1_Y, Y => AND2_24_Y);
    
    XNOR2_0 : XNOR2
      port map(A => MEM_RADDR_0_net, B => WBINNXTSHIFT_0_net, Y
         => XNOR2_0_Y);
    
    DFN1E1C0_Q_39_inst : DFN1E1C0
      port map(D => QXI_39_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_5, E => DVLDI_1, Q => 
        \Z\\Fifo_wr_0_Q_[39]\\\);
    
    AND2_31 : AND2
      port map(A => WBINNXTSHIFT_2_net, B => INV_4_Y, Y => 
        AND2_31_Y);
    
    GND_i : GND
      port map(Y => \GND\);
    
    XOR2_WBINNXTSHIFT_0_inst : XOR2
      port map(A => MEM_WADDR_0_net, B => MEMORYWE, Y => 
        WBINNXTSHIFT_0_net);
    
    XOR2_18 : XOR2
      port map(A => MEM_WADDR_1_net, B => Fifo_rd_GND, Y => 
        XOR2_18_Y);
    
    DFN1E1C0_Q_41_inst : DFN1E1C0
      port map(D => QXI_41_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_6, E => DVLDI_1, Q => 
        \Z\\Fifo_wr_0_Q_[41]\\\);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    NAND3A_0 : NAND3A
      port map(A => WDIFF_1_net, B => Fifo_rd_GND, C => OR2A_1_Y, 
        Y => NAND3A_0_Y);
    
    DFN1E1C0_Q_45_inst : DFN1E1C0
      port map(D => QXI_45_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_6, E => DVLDI_1, Q => 
        \Z\\Fifo_wr_0_Q_[45]\\\);
    
    XOR2_RBINNXTSHIFT_2_inst : XOR2
      port map(A => XOR2_10_Y, B => AO1_8_Y, Y => 
        RBINNXTSHIFT_2_net);
    
    DFN1E1C0_Q_67_inst : DFN1E1C0
      port map(D => QXI_67_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n, E => DVLDI_2, Q => 
        \Z\\Fifo_wr_0_Q_[67]\\\);
    
    MEMREBUBBLE : INV
      port map(A => MEMORYRE, Y => MEMRENEG);
    
    DFN1E1C0_Q_20_inst : DFN1E1C0
      port map(D => QXI_20_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_5, E => DVLDI_0, Q => 
        \Z\\Fifo_wr_0_Q_[20]\\\);
    
    DFN1E1C0_Q_63_inst : DFN1E1C0
      port map(D => QXI_63_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n, E => DVLDI_2, Q => 
        \Z\\Fifo_wr_0_Q_[63]\\\);
    
    XOR2_RBINNXTSHIFT_0_inst : XOR2
      port map(A => MEM_RADDR_0_net, B => MEMORYRE, Y => 
        RBINNXTSHIFT_0_net);
    
    XOR2_WBINNXTSHIFT_1_inst : XOR2
      port map(A => XOR2_0_Y, B => AND2_8_Y, Y => 
        WBINNXTSHIFT_1_net);
    
    DFN1E1C0_Q_30_inst : DFN1E1C0
      port map(D => QXI_30_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_5, E => DVLDI_0, Q => 
        \Z\\Fifo_wr_0_Q_[30]\\\);
    
    AND2_3 : AND2
      port map(A => MEM_WADDR_2_net, B => Fifo_rd_GND, Y => 
        AND2_3_Y);
    
    DFN1E1C0_Q_28_inst : DFN1E1C0
      port map(D => QXI_28_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_5, E => DVLDI_0, Q => 
        \Z\\Fifo_wr_0_Q_[28]\\\);
    
    DFN1E1C0_Q_46_inst : DFN1E1C0
      port map(D => QXI_46_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_6, E => DVLDI_1, Q => 
        \Z\\Fifo_wr_0_Q_[46]\\\);
    
    XNOR2_6 : XNOR2
      port map(A => RBINNXTSHIFT_3_net, B => MEM_WADDR_3_net, Y
         => XNOR2_6_Y);
    
    OA1C_0 : OA1C
      port map(A => Fifo_rd_VCC, B => WDIFF_3_net, C => 
        Fifo_rd_GND, Y => OA1C_0_Y);
    
    INV_4 : INV
      port map(A => MEM_RADDR_2_net, Y => INV_4_Y);
    
    OR2A_1 : OR2A
      port map(A => WDIFF_2_net, B => Fifo_rd_GND, Y => OR2A_1_Y);
    
    DFN1E1C0_Q_38_inst : DFN1E1C0
      port map(D => QXI_38_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_5, E => DVLDI_1, Q => 
        \Z\\Fifo_wr_0_Q_[38]\\\);
    
    DFN1E1C0_Q_42_inst : DFN1E1C0
      port map(D => QXI_42_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_6, E => DVLDI_1, Q => 
        \Z\\Fifo_wr_0_Q_[42]\\\);
    
    DFN1E1C0_Q_51_inst : DFN1E1C0
      port map(D => QXI_51_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_6, E => DVLDI_1, Q => 
        \Z\\Fifo_wr_0_Q_[51]\\\);
    
    XOR2_9 : XOR2
      port map(A => WBINNXTSHIFT_3_net, B => INV_2_Y, Y => 
        XOR2_9_Y);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    XOR2_RBINNXTSHIFT_1_inst : XOR2
      port map(A => XOR2_29_Y, B => AND2_28_Y, Y => 
        RBINNXTSHIFT_1_net);
    
    XNOR2_4 : XNOR2
      port map(A => Fifo_rd_VCC, B => WDIFF_3_net, Y => XNOR2_4_Y);
    
    DFN1E1C0_Q_55_inst : DFN1E1C0
      port map(D => QXI_55_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_6, E => DVLDI_2, Q => 
        \Z\\Fifo_wr_0_Q_[55]\\\);
    
    DFN1E1C0_Q_1_inst : DFN1E1C0
      port map(D => QXI_1_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_4, E => DVLDI_0, Q => 
        \Z\\Fifo_wr_0_Q_[1]\\\);
    
    DFN1C0_MEM_WADDR_4_inst : DFN1C0
      port map(D => WBINNXTSHIFT_4_net, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => 
        Main_ctl4SD_0_fifo_rst_n_4, Q => MEM_WADDR_4_net);
    
    DFN1E1C0_Q_4_inst : DFN1E1C0
      port map(D => QXI_4_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_6, E => DVLDI_1, Q => 
        \Z\\Fifo_wr_0_Q_[4]\\\);
    
    XOR2_13 : XOR2
      port map(A => MEM_WADDR_2_net, B => Fifo_rd_GND, Y => 
        XOR2_13_Y);
    
    DFN1E1C0_Q_8_inst : DFN1E1C0
      port map(D => QXI_8_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n, E => DVLDI_2, Q => 
        \Z\\Fifo_wr_0_Q_[8]\\\);
    
    XOR2_WBINNXTSHIFT_3_inst : XOR2
      port map(A => XOR2_32_Y, B => AO1_4_Y, Y => 
        WBINNXTSHIFT_3_net);
    
    XOR2_WDIFF_4_inst : XOR2
      port map(A => XOR2_21_Y, B => AO1_6_Y, Y => WDIFF_4_net);
    
    DFN1E1C0_Q_56_inst : DFN1E1C0
      port map(D => QXI_56_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_6, E => DVLDI_2, Q => 
        \Z\\Fifo_wr_0_Q_[56]\\\);
    
    AO1_3 : AO1
      port map(A => AND2_12_Y, B => AO1_0_Y, C => AO1_10_Y, Y => 
        AO1_3_Y);
    
    DFN1E1C0_Q_70_inst : DFN1E1C0
      port map(D => QXI_70_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n, E => DVLDI_2, Q => 
        \Z\\Fifo_wr_0_Q_[70]\\\);
    
    DFN1E1C0_Q_47_inst : DFN1E1C0
      port map(D => QXI_47_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_6, E => DVLDI_1, Q => 
        \Z\\Fifo_wr_0_Q_[47]\\\);
    
    DFN1E1C0_Q_52_inst : DFN1E1C0
      port map(D => QXI_52_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_6, E => DVLDI_1, Q => 
        \Z\\Fifo_wr_0_Q_[52]\\\);
    
    AO1C_0 : AO1C
      port map(A => Fifo_rd_GND, B => WDIFF_1_net, C => 
        Fifo_rd_GND, Y => AO1C_0_Y);
    
    DFN1E1C0_Q_7_inst : DFN1E1C0
      port map(D => QXI_7_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n, E => DVLDI_2, Q => 
        \Z\\Fifo_wr_0_Q_[7]\\\);
    
    DFN1E1C0_Q_43_inst : DFN1E1C0
      port map(D => QXI_43_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_6, E => DVLDI_1, Q => 
        \Z\\Fifo_wr_0_Q_[43]\\\);
    
    AND2_13 : AND2
      port map(A => MEM_RADDR_1_net, B => Fifo_rd_GND, Y => 
        AND2_13_Y);
    
    DFN1E1C0_Q_11_inst : DFN1E1C0
      port map(D => QXI_11_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_4, E => DVLDI_0, Q => 
        \Z\\Fifo_wr_0_Q_[11]\\\);
    
    XOR2_10 : XOR2
      port map(A => MEM_RADDR_2_net, B => Fifo_rd_GND, Y => 
        XOR2_10_Y);
    
    XNOR2_1 : XNOR2
      port map(A => Fifo_rd_GND, B => WDIFF_4_net, Y => XNOR2_1_Y);
    
    XOR2_RBINNXTSHIFT_3_inst : XOR2
      port map(A => XOR2_28_Y, B => AO1_13_Y, Y => 
        RBINNXTSHIFT_3_net);
    
    DFN1E1C0_Q_15_inst : DFN1E1C0
      port map(D => QXI_15_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_4, E => DVLDI_0, Q => 
        \Z\\Fifo_wr_0_Q_[15]\\\);
    
    DFN1E1C0_Q_69_inst : DFN1E1C0
      port map(D => QXI_69_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n, E => DVLDI_2, Q => 
        \Z\\Fifo_wr_0_Q_[69]\\\);
    
    AND2_MEMORYRE : AND2
      port map(A => NAND2_1_Y, B => Sdram_cmd_0_WFifo_re, Y => 
        MEMORYRE);
    
    XOR2_7 : XOR2
      port map(A => WBINNXTSHIFT_2_net, B => INV_4_Y, Y => 
        XOR2_7_Y);
    
    XOR2_14 : XOR2
      port map(A => WBINNXTSHIFT_1_net, B => INV_1_Y, Y => 
        XOR2_14_Y);
    
    XOR2_11 : XOR2
      port map(A => MEM_WADDR_2_net, B => Fifo_rd_GND, Y => 
        XOR2_11_Y);
    
    XNOR2_3 : XNOR2
      port map(A => RBINNXTSHIFT_0_net, B => MEM_WADDR_0_net, Y
         => XNOR2_3_Y);
    
    DFN1E1C0_Q_24_inst : DFN1E1C0
      port map(D => QXI_24_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_5, E => DVLDI_0, Q => 
        \Z\\Fifo_wr_0_Q_[24]\\\);
    
    DFN1E1C0_Q_34_inst : DFN1E1C0
      port map(D => QXI_34_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_5, E => DVLDI_1, Q => 
        \Z\\Fifo_wr_0_Q_[34]\\\);
    
    DFN1E1C0_Q_57_inst : DFN1E1C0
      port map(D => QXI_57_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_6, E => DVLDI_2, Q => 
        \Z\\Fifo_wr_0_Q_[57]\\\);
    
    DFN1E1C0_Q_16_inst : DFN1E1C0
      port map(D => QXI_16_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_4, E => DVLDI_0, Q => 
        \Z\\Fifo_wr_0_Q_[16]\\\);
    
    DFN1C0_MEM_RADDR_3_inst : DFN1C0
      port map(D => RBINNXTSHIFT_3_net, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => 
        Main_ctl4SD_0_fifo_rst_n_4, Q => MEM_RADDR_3_net);
    
    AO1_6 : AO1
      port map(A => XOR2_3_Y, B => AO1_7_Y, C => AND2_9_Y, Y => 
        AO1_6_Y);
    
    DFN1E1C0_Q_12_inst : DFN1E1C0
      port map(D => QXI_12_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_4, E => DVLDI_0, Q => 
        \Z\\Fifo_wr_0_Q_[12]\\\);
    
    DFN1E1C0_Q_53_inst : DFN1E1C0
      port map(D => QXI_53_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_6, E => DVLDI_2, Q => 
        \Z\\Fifo_wr_0_Q_[53]\\\);
    
    XOR2_WBINNXTSHIFT_4_inst : XOR2
      port map(A => XOR2_16_Y, B => AO1_3_Y, Y => 
        WBINNXTSHIFT_4_net);
    
    DFN1E1C0_Q_60_inst : DFN1E1C0
      port map(D => QXI_60_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_6, E => DVLDI_2, Q => 
        \Z\\Fifo_wr_0_Q_[60]\\\);
    
    XOR2_32 : XOR2
      port map(A => MEM_WADDR_3_net, B => Fifo_rd_GND, Y => 
        XOR2_32_Y);
    
    OR3_0 : OR3
      port map(A => AND2_22_Y, B => AND2_17_Y, C => AND2_2_Y, Y
         => OR3_0_Y);
    
    AND2_9 : AND2
      port map(A => WBINNXTSHIFT_3_net, B => INV_2_Y, Y => 
        AND2_9_Y);
    
    RAM512X18_QXI_71_inst : RAM512X18
      port map(RADDR8 => Fifo_rd_GND, RADDR7 => Fifo_rd_GND, 
        RADDR6 => Fifo_rd_GND, RADDR5 => Fifo_rd_GND, RADDR4 => 
        Fifo_rd_GND, RADDR3 => MEM_RADDR_3_net, RADDR2 => 
        MEM_RADDR_2_net, RADDR1 => MEM_RADDR_1_net, RADDR0 => 
        MEM_RADDR_0_net, WADDR8 => Fifo_rd_GND, WADDR7 => 
        Fifo_rd_GND, WADDR6 => Fifo_rd_GND, WADDR5 => Fifo_rd_GND, 
        WADDR4 => Fifo_rd_GND, WADDR3 => MEM_WADDR_3_net, WADDR2
         => MEM_WADDR_2_net, WADDR1 => MEM_WADDR_1_net, WADDR0
         => MEM_WADDR_0_net, WD17 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[71]\\\, WD16 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[70]\\\, WD15 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[69]\\\, WD14 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[68]\\\, WD13 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[67]\\\, WD12 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[66]\\\, WD11 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[65]\\\, WD10 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[64]\\\, WD9 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[63]\\\, WD8 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[62]\\\, WD7 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[61]\\\, WD6 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[60]\\\, WD5 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[59]\\\, WD4 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[58]\\\, WD3 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[57]\\\, WD2 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[56]\\\, WD1 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[55]\\\, WD0 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[54]\\\, RW0 => Fifo_rd_GND, 
        RW1 => Fifo_rd_VCC, WW0 => Fifo_rd_GND, WW1 => 
        Fifo_rd_VCC, PIPE => Fifo_rd_GND, REN => MEMRENEG, WEN
         => MEMWENEG, RCLK => PLL_Test1_0_Sys_66M_Clk, WCLK => 
        PLL_Test1_0_Sys_66M_Clk, RESET => 
        Main_ctl4SD_0_fifo_rst_n, RD17 => QXI_71_net, RD16 => 
        QXI_70_net, RD15 => QXI_69_net, RD14 => QXI_68_net, RD13
         => QXI_67_net, RD12 => QXI_66_net, RD11 => QXI_65_net, 
        RD10 => QXI_64_net, RD9 => QXI_63_net, RD8 => QXI_62_net, 
        RD7 => QXI_61_net, RD6 => QXI_60_net, RD5 => QXI_59_net, 
        RD4 => QXI_58_net, RD3 => QXI_57_net, RD2 => QXI_56_net, 
        RD1 => QXI_55_net, RD0 => QXI_54_net);
    
    NOR3A_0 : NOR3A
      port map(A => OR2A_1_Y, B => AO1C_0_Y, C => WDIFF_0_net, Y
         => NOR3A_0_Y);
    
    DFN1E1C0_Q_68_inst : DFN1E1C0
      port map(D => QXI_68_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n, E => DVLDI_2, Q => 
        \Z\\Fifo_wr_0_Q_[68]\\\);
    
    DFN1C0_AFULL : DFN1C0
      port map(D => OR2_0_Y, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => Main_ctl4SD_0_fifo_rst_n_3, Q => Fifo_wr_0_AFULL);
    
    INV_2 : INV
      port map(A => MEM_RADDR_3_net, Y => INV_2_Y);
    
    DFN1C0_MEM_WADDR_1_inst : DFN1C0
      port map(D => WBINNXTSHIFT_1_net, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => 
        Main_ctl4SD_0_fifo_rst_n_4, Q => MEM_WADDR_1_net);
    
    NAND3A_1 : NAND3A
      port map(A => NOR3A_0_Y, B => OR2A_0_Y, C => NAND3A_0_Y, Y
         => NAND3A_1_Y);
    
    NAND2_0 : NAND2
      port map(A => DFN1C0_FULL_1, B => Fifo_rd_VCC, Y => 
        NAND2_0_Y);
    
    DFN1E1C0_Q_3_inst : DFN1E1C0
      port map(D => QXI_3_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_5, E => DVLDI_1, Q => 
        \Z\\Fifo_wr_0_Q_[3]\\\);
    
    XOR2_RBINNXTSHIFT_4_inst : XOR2
      port map(A => XOR2_36_Y, B => AO1_5_Y, Y => 
        RBINNXTSHIFT_4_net);
    
    DFN1C0_DVLDI : DFN1C0
      port map(D => AND2A_1_Y, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_3, Q => DVLDI);
    
    XNOR2_10 : XNOR2
      port map(A => RBINNXTSHIFT_4_net, B => MEM_WADDR_4_net, Y
         => XNOR2_10_Y);
    
    AND2_MEMORYWE : AND2
      port map(A => NAND2_0_Y, B => Main_ctl4SD_0_Fifo_wr, Y => 
        MEMORYWE);
    
    DFN1E1C0_Q_49_inst : DFN1E1C0
      port map(D => QXI_49_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_6, E => DVLDI_1, Q => 
        \Z\\Fifo_wr_0_Q_[49]\\\);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    DFN1E1C0_Q_17_inst : DFN1E1C0
      port map(D => QXI_17_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_4, E => DVLDI_0, Q => 
        \Z\\Fifo_wr_0_Q_[17]\\\);
    
    AO1_0 : AO1
      port map(A => XOR2_18_Y, B => AND2_8_Y, C => AND2_18_Y, Y
         => AO1_0_Y);
    
    XOR2_29 : XOR2
      port map(A => MEM_RADDR_1_net, B => Fifo_rd_GND, Y => 
        XOR2_29_Y);
    
    XOR2_2 : XOR2
      port map(A => MEM_RADDR_1_net, B => Fifo_rd_GND, Y => 
        XOR2_2_Y);
    
    DFN1C0_MEM_WADDR_0_inst : DFN1C0
      port map(D => WBINNXTSHIFT_0_net, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => 
        Main_ctl4SD_0_fifo_rst_n_4, Q => MEM_WADDR_0_net);
    
    DFN1E1C0_Q_13_inst : DFN1E1C0
      port map(D => QXI_13_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_4, E => DVLDI_0, Q => 
        \Z\\Fifo_wr_0_Q_[13]\\\);
    
    AND2A_0 : AND2A
      port map(A => Fifo_rd_GND, B => WDIFF_4_net, Y => AND2A_0_Y);
    
    OA1A_0 : OA1A
      port map(A => Fifo_rd_VCC, B => WDIFF_3_net, C => 
        WDIFF_4_net, Y => OA1A_0_Y);
    
    AOI1_0 : AOI1
      port map(A => AND2_6_Y, B => NAND3A_1_Y, C => NOR3_0_Y, Y
         => AOI1_0_Y);
    
    AO1_10 : AO1
      port map(A => XOR2_35_Y, B => AND2_3_Y, C => AND2_1_Y, Y
         => AO1_10_Y);
    
    XOR2_35 : XOR2
      port map(A => MEM_WADDR_3_net, B => Fifo_rd_GND, Y => 
        XOR2_35_Y);
    
    DFN1P0_EMPTY : DFN1P0
      port map(D => EMPTYINT, CLK => PLL_Test1_0_Sys_66M_Clk, PRE
         => Main_ctl4SD_0_fifo_rst_n, Q => DFN1P0_EMPTY_1);
    
    AND2_17 : AND2
      port map(A => WBINNXTSHIFT_1_net, B => INV_3_Y, Y => 
        AND2_17_Y);
    
    DFN1E1C0_Q_40_inst : DFN1E1C0
      port map(D => QXI_40_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_5, E => DVLDI_1, Q => 
        \Z\\Fifo_wr_0_Q_[40]\\\);
    
    NOR2A_0 : NOR2A
      port map(A => MEM_RADDR_0_net, B => WBINNXTSHIFT_0_net, Y
         => NOR2A_0_Y);
    
    AO1_13 : AO1
      port map(A => XOR2_4_Y, B => AO1_8_Y, C => AND2_4_Y, Y => 
        AO1_13_Y);
    
    DFN1C0_MEM_WADDR_3_inst : DFN1C0
      port map(D => WBINNXTSHIFT_3_net, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => 
        Main_ctl4SD_0_fifo_rst_n_4, Q => MEM_WADDR_3_net);
    
    DFN1E1C0_Q_48_inst : DFN1E1C0
      port map(D => QXI_48_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_6, E => DVLDI_1, Q => 
        \Z\\Fifo_wr_0_Q_[48]\\\);
    
    DFN1E1C0_Q_9_inst : DFN1E1C0
      port map(D => QXI_9_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n, E => DVLDI_2, Q => 
        \Z\\Fifo_wr_0_Q_[9]\\\);
    
    DFN1E1C0_Q_59_inst : DFN1E1C0
      port map(D => QXI_59_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_6, E => DVLDI_2, Q => 
        \Z\\Fifo_wr_0_Q_[59]\\\);
    
    XNOR2_WDIFF_1_inst : XNOR2
      port map(A => XOR2_14_Y, B => NOR2A_0_Y, Y => WDIFF_1_net);
    
    OR2A_0 : OR2A
      port map(A => Fifo_rd_GND, B => WDIFF_2_net, Y => OR2A_0_Y);
    
    XNOR2_7 : XNOR2
      port map(A => MEM_RADDR_1_net, B => WBINNXTSHIFT_1_net, Y
         => XNOR2_7_Y);
    
    DFN1C0_DVLDI_RNI1QG2 : BUFF
      port map(A => DVLDI, Y => DVLDI_1);
    
    DFN1E1C0_Q_64_inst : DFN1E1C0
      port map(D => QXI_64_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n, E => DVLDI_2, Q => 
        \Z\\Fifo_wr_0_Q_[64]\\\);
    
    DFN1C0_MEM_RADDR_2_inst : DFN1C0
      port map(D => RBINNXTSHIFT_2_net, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => 
        Main_ctl4SD_0_fifo_rst_n_4, Q => MEM_RADDR_2_net);
    
    AND2_4 : AND2
      port map(A => MEM_RADDR_2_net, B => Fifo_rd_GND, Y => 
        AND2_4_Y);
    
    AND2_FULLINT : AND2
      port map(A => AND2_7_Y, B => XOR2_23_Y, Y => FULLINT);
    
    DFN1C0_MEM_RADDR_1_inst : DFN1C0
      port map(D => RBINNXTSHIFT_1_net, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => 
        Main_ctl4SD_0_fifo_rst_n_4, Q => MEM_RADDR_1_net);
    
    XNOR2_5 : XNOR2
      port map(A => RBINNXTSHIFT_2_net, B => MEM_WADDR_2_net, Y
         => XNOR2_5_Y);
    
    DFN1E1C0_Q_21_inst : DFN1E1C0
      port map(D => QXI_21_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_5, E => DVLDI_0, Q => 
        \Z\\Fifo_wr_0_Q_[21]\\\);
    
    AO1_5 : AO1
      port map(A => AND2_24_Y, B => AO1_8_Y, C => AO1_11_Y, Y => 
        AO1_5_Y);
    
    DFN1E1C0_Q_50_inst : DFN1E1C0
      port map(D => QXI_50_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_6, E => DVLDI_1, Q => 
        \Z\\Fifo_wr_0_Q_[50]\\\);
    
    AND2_8 : AND2
      port map(A => MEM_WADDR_0_net, B => MEMORYWE, Y => AND2_8_Y);
    
    XOR2_3 : XOR2
      port map(A => WBINNXTSHIFT_3_net, B => INV_2_Y, Y => 
        XOR2_3_Y);
    
    RAM512X18_QXI_35_inst : RAM512X18
      port map(RADDR8 => Fifo_rd_GND, RADDR7 => Fifo_rd_GND, 
        RADDR6 => Fifo_rd_GND, RADDR5 => Fifo_rd_GND, RADDR4 => 
        Fifo_rd_GND, RADDR3 => MEM_RADDR_3_net, RADDR2 => 
        MEM_RADDR_2_net, RADDR1 => MEM_RADDR_1_net, RADDR0 => 
        MEM_RADDR_0_net, WADDR8 => Fifo_rd_GND, WADDR7 => 
        Fifo_rd_GND, WADDR6 => Fifo_rd_GND, WADDR5 => Fifo_rd_GND, 
        WADDR4 => Fifo_rd_GND, WADDR3 => MEM_WADDR_3_net, WADDR2
         => MEM_WADDR_2_net, WADDR1 => MEM_WADDR_1_net, WADDR0
         => MEM_WADDR_0_net, WD17 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[35]\\\, WD16 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[34]\\\, WD15 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[33]\\\, WD14 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[32]\\\, WD13 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[31]\\\, WD12 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[30]\\\, WD11 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[29]\\\, WD10 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[28]\\\, WD9 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[27]\\\, WD8 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[26]\\\, WD7 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[25]\\\, WD6 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[24]\\\, WD5 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[23]\\\, WD4 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[22]\\\, WD3 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[21]\\\, WD2 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[20]\\\, WD1 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[19]\\\, WD0 => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[18]\\\, RW0 => Fifo_rd_GND, 
        RW1 => Fifo_rd_VCC, WW0 => Fifo_rd_GND, WW1 => 
        Fifo_rd_VCC, PIPE => Fifo_rd_GND, REN => MEMRENEG, WEN
         => MEMWENEG, RCLK => PLL_Test1_0_Sys_66M_Clk, WCLK => 
        PLL_Test1_0_Sys_66M_Clk, RESET => 
        Main_ctl4SD_0_fifo_rst_n, RD17 => QXI_35_net, RD16 => 
        QXI_34_net, RD15 => QXI_33_net, RD14 => QXI_32_net, RD13
         => QXI_31_net, RD12 => QXI_30_net, RD11 => QXI_29_net, 
        RD10 => QXI_28_net, RD9 => QXI_27_net, RD8 => QXI_26_net, 
        RD7 => QXI_25_net, RD6 => QXI_24_net, RD5 => QXI_23_net, 
        RD4 => QXI_22_net, RD3 => QXI_21_net, RD2 => QXI_20_net, 
        RD1 => QXI_19_net, RD0 => QXI_18_net);
    
    DFN1E1C0_Q_31_inst : DFN1E1C0
      port map(D => QXI_31_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_5, E => DVLDI_1, Q => 
        \Z\\Fifo_wr_0_Q_[31]\\\);
    
    DFN1E1C0_Q_25_inst : DFN1E1C0
      port map(D => QXI_25_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_5, E => DVLDI_0, Q => 
        \Z\\Fifo_wr_0_Q_[25]\\\);
    
    DFN1E1C0_Q_58_inst : DFN1E1C0
      port map(D => QXI_58_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_6, E => DVLDI_2, Q => 
        \Z\\Fifo_wr_0_Q_[58]\\\);
    
    DFN1E1C0_Q_35_inst : DFN1E1C0
      port map(D => QXI_35_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_5, E => DVLDI_1, Q => 
        \Z\\Fifo_wr_0_Q_[35]\\\);
    
    DFN1E1C0_Q_19_inst : DFN1E1C0
      port map(D => QXI_19_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_4, E => DVLDI_0, Q => 
        \Z\\Fifo_wr_0_Q_[19]\\\);
    
    XOR2_28 : XOR2
      port map(A => MEM_RADDR_3_net, B => Fifo_rd_GND, Y => 
        XOR2_28_Y);
    
    XOR2_WDIFF_2_inst : XOR2
      port map(A => XOR2_20_Y, B => OR3_0_Y, Y => WDIFF_2_net);
    
    DFN1E1C0_Q_26_inst : DFN1E1C0
      port map(D => QXI_26_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_5, E => DVLDI_0, Q => 
        \Z\\Fifo_wr_0_Q_[26]\\\);
    
    DFN1E1C0_Q_22_inst : DFN1E1C0
      port map(D => QXI_22_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_5, E => DVLDI_0, Q => 
        \Z\\Fifo_wr_0_Q_[22]\\\);
    
    DFN1E1C0_Q_36_inst : DFN1E1C0
      port map(D => QXI_36_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_5, E => DVLDI_1, Q => 
        \Z\\Fifo_wr_0_Q_[36]\\\);
    
    AND2_21 : AND2
      port map(A => MEM_RADDR_3_net, B => Fifo_rd_GND, Y => 
        AND2_21_Y);
    
    XOR2_WDIFF_3_inst : XOR2
      port map(A => XOR2_9_Y, B => AO1_7_Y, Y => WDIFF_3_net);
    
    DFN1E1C0_Q_32_inst : DFN1E1C0
      port map(D => QXI_32_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_5, E => DVLDI_1, Q => 
        \Z\\Fifo_wr_0_Q_[32]\\\);
    
    DFN1E1C0_Q_6_inst : DFN1E1C0
      port map(D => QXI_6_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n, E => DVLDI_2, Q => 
        \Z\\Fifo_wr_0_Q_[6]\\\);
    
    XOR2_0 : XOR2
      port map(A => MEM_WADDR_1_net, B => Fifo_rd_GND, Y => 
        XOR2_0_Y);
    
    NAND2_1 : NAND2
      port map(A => DFN1P0_EMPTY_1, B => Fifo_rd_VCC, Y => 
        NAND2_1_Y);
    
    DFN1E1C0_Q_44_inst : DFN1E1C0
      port map(D => QXI_44_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_6, E => DVLDI_1, Q => 
        \Z\\Fifo_wr_0_Q_[44]\\\);
    
    DFN1C0_MEM_RADDR_4_inst : DFN1C0
      port map(D => RBINNXTSHIFT_4_net, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => 
        Main_ctl4SD_0_fifo_rst_n_4, Q => MEM_RADDR_4_net);
    
    DFN1E1C0_Q_10_inst : DFN1E1C0
      port map(D => QXI_10_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_4, E => DVLDI_0, Q => 
        \Z\\Fifo_wr_0_Q_[10]\\\);
    
    AO1_4 : AO1
      port map(A => XOR2_11_Y, B => AO1_0_Y, C => AND2_3_Y, Y => 
        AO1_4_Y);
    
    DFN1E1C0_Q_71_inst : DFN1E1C0
      port map(D => QXI_71_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n, E => DVLDI_2, Q => 
        \Z\\Fifo_wr_0_Q_[71]\\\);
    
    DFN1E1C0_Q_18_inst : DFN1E1C0
      port map(D => QXI_18_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_4, E => DVLDI_0, Q => 
        \Z\\Fifo_wr_0_Q_[18]\\\);
    
    XOR2_36 : XOR2
      port map(A => MEM_RADDR_4_net, B => Fifo_rd_GND, Y => 
        XOR2_36_Y);
    
    XNOR2_8 : XNOR2
      port map(A => MEM_RADDR_3_net, B => WBINNXTSHIFT_3_net, Y
         => XNOR2_8_Y);
    
    XOR2_WDIFF_0_inst : XOR2
      port map(A => WBINNXTSHIFT_0_net, B => MEM_RADDR_0_net, Y
         => WDIFF_0_net);
    
    AND2_28 : AND2
      port map(A => MEM_RADDR_0_net, B => MEMORYRE, Y => 
        AND2_28_Y);
    
    AND2_25 : AND2
      port map(A => AND3_1_Y, B => XNOR2_6_Y, Y => AND2_25_Y);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3;
use proasic3.all;

entity WaveGenSingleZ6 is

    port( PrState_3               : in    std_logic;
          Clock_Y_c               : out   std_logic;
          PLL_Test1_0_SysRst_O    : in    std_logic;
          PLL_Test1_0_Sys_66M_Clk : in    std_logic;
          RowReadOutEn            : in    std_logic;
          RowReadOutEn_0          : in    std_logic
        );

end WaveGenSingleZ6;

architecture DEF_ARCH of WaveGenSingleZ6 is 

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \PrState_ns_tz_0[2]\, \DelayCnt_RNIEUP7[0]_net_1\, 
        \Phase1Cnt_RNI6GC8[0]_net_1\, \PrState_RNO_0[1]_net_1\, 
        N_84, N_85, \PrState_ns[2]\, \PrState_ns_a3_1_0[2]\, N_73, 
        \CycCnt[0]_net_1\, N_75, \PrState[3]_net_1\, 
        \DelayCnt[0]_net_1\, \PrState[1]_net_1\, 
        \Phase2Cnt[0]_net_1\, \CycCnt_RNO_0[0]\, 
        \PrState_RNO_1[3]\, \PrState[2]_net_1\, 
        \Phase1Cnt[0]_net_1\, \GND\, \VCC\, GND_0, VCC_0
         : std_logic;

begin 


    \DelayCnt_RNIEUP7[0]\ : NOR2A
      port map(A => \PrState[3]_net_1\, B => \DelayCnt[0]_net_1\, 
        Y => \DelayCnt_RNIEUP7[0]_net_1\);
    
    \PrState_RNO[2]\ : OA1
      port map(A => \PrState_ns_a3_1_0[2]\, B => 
        \PrState_ns_tz_0[2]\, C => RowReadOutEn_0, Y => 
        \PrState_ns[2]\);
    
    \DelayCnt[0]\ : DFN1C0
      port map(D => \DelayCnt_RNIEUP7[0]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \DelayCnt[0]_net_1\);
    
    WFO : DFN1C0
      port map(D => \PrState[2]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => Clock_Y_c);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    \PrState[3]\ : DFN1C0
      port map(D => \PrState_RNO_1[3]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \PrState[3]_net_1\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \PrState[1]\ : DFN1C0
      port map(D => \PrState_RNO_0[1]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \PrState[1]_net_1\);
    
    \PrState_RNO_1[1]\ : NOR2
      port map(A => \PrState[1]_net_1\, B => \Phase1Cnt[0]_net_1\, 
        Y => N_85);
    
    \PrState_RNO_0[1]\ : AOI1
      port map(A => \PrState[1]_net_1\, B => \Phase2Cnt[0]_net_1\, 
        C => \PrState[2]_net_1\, Y => N_84);
    
    \CycCnt[0]\ : DFN1C0
      port map(D => \CycCnt_RNO_0[0]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \CycCnt[0]_net_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \PrState_RNO[1]\ : NOR3A
      port map(A => RowReadOutEn_0, B => N_84, C => N_85, Y => 
        \PrState_RNO_0[1]_net_1\);
    
    \PrState_RNO[3]\ : OA1
      port map(A => N_75, B => PrState_3, C => RowReadOutEn, Y
         => \PrState_RNO_1[3]\);
    
    \CycCnt_RNO[0]\ : XA1B
      port map(A => \CycCnt[0]_net_1\, B => N_73, C => PrState_3, 
        Y => \CycCnt_RNO_0[0]\);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    \Phase1Cnt_RNI6GC8[0]\ : NOR2A
      port map(A => \PrState[2]_net_1\, B => \Phase1Cnt[0]_net_1\, 
        Y => \Phase1Cnt_RNI6GC8[0]_net_1\);
    
    \PrState_RNO_1[2]\ : OR2
      port map(A => \DelayCnt_RNIEUP7[0]_net_1\, B => 
        \Phase1Cnt_RNI6GC8[0]_net_1\, Y => \PrState_ns_tz_0[2]\);
    
    \Phase1Cnt[0]\ : DFN1C0
      port map(D => \Phase1Cnt_RNI6GC8[0]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \Phase1Cnt[0]_net_1\);
    
    \Phase2Cnt[0]\ : DFN1C0
      port map(D => N_73, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase2Cnt[0]_net_1\);
    
    \PrState_RNO_0[2]\ : NOR2B
      port map(A => N_73, B => \CycCnt[0]_net_1\, Y => 
        \PrState_ns_a3_1_0[2]\);
    
    \Phase2Cnt_RNI05E8[0]\ : NOR2A
      port map(A => \PrState[1]_net_1\, B => \Phase2Cnt[0]_net_1\, 
        Y => N_73);
    
    \PrState_RNO_0[3]\ : NOR2B
      port map(A => \PrState[3]_net_1\, B => \DelayCnt[0]_net_1\, 
        Y => N_75);
    
    \PrState[2]\ : DFN1C0
      port map(D => \PrState_ns[2]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \PrState[2]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3;
use proasic3.all;

entity sampleEn_dly is

    port( sampleEn_dly_VCC        : in    std_logic;
          sampleEn_dly_GND        : in    std_logic;
          AdcCLkEn                : in    std_logic;
          PLL_Test1_0_ADC_66M_Clk : in    std_logic;
          DRY_c_c                 : out   std_logic
        );

end sampleEn_dly;

architecture DEF_ARCH of sampleEn_dly is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CLKDLY
    port( CLK    : in    std_logic := 'U';
          GL     : out   std_logic;
          DLYGL0 : in    std_logic := 'U';
          DLYGL1 : in    std_logic := 'U';
          DLYGL2 : in    std_logic := 'U';
          DLYGL3 : in    std_logic := 'U';
          DLYGL4 : in    std_logic := 'U'
        );
  end component;

    signal AdcCLKEn_DLY, \GND\, \VCC\, GND_0, VCC_0 : std_logic;

begin 


    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    Inst1_RNIBMI8 : NOR2B
      port map(A => PLL_Test1_0_ADC_66M_Clk, B => AdcCLKEn_DLY, Y
         => DRY_c_c);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    Inst1 : CLKDLY
      port map(CLK => AdcCLkEn, GL => AdcCLKEn_DLY, DLYGL0 => 
        sampleEn_dly_GND, DLYGL1 => sampleEn_dly_GND, DLYGL2 => 
        sampleEn_dly_GND, DLYGL3 => sampleEn_dly_VCC, DLYGL4 => 
        sampleEn_dly_GND);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3;
use proasic3.all;

entity WaveGenSingleZ0 is

    port( PrState_4               : out   std_logic;
          PrState_0               : out   std_logic_vector(4 to 4);
          Adc_RdEn_inter          : out   std_logic;
          RowReadOutEn            : in    std_logic;
          RowReadOutEn_0          : in    std_logic;
          PLL_Test1_0_SysRst_O    : in    std_logic;
          RowReadOutEn_i          : in    std_logic;
          PLL_Test1_0_Sys_66M_Clk : in    std_logic
        );

end WaveGenSingleZ0;

architecture DEF_ARCH of WaveGenSingleZ0 is 

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component AX1E
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \PrState_ns_0_i_a2_0_0_0[1]\, \DelayCnt[4]_net_1\, 
        \DelayCnt[2]_net_1\, \DelayCnt[3]_net_1\, 
        \CycCnt_5_i_o2_0[0]\, \PrState[0]_net_1\, 
        \Phase2Cnt[0]_net_1\, N_68, \PrState[1]_net_1\, N_10, 
        N_63, N_64, N_50, \PrState_0[4]_net_1\, N_58, 
        \PrState[3]_net_1\, \PrState[2]_net_1\, N_36, N_48, 
        \Phase1Cnt[8]_net_1\, N_34, N_47, \Phase1Cnt[7]_net_1\, 
        N_32, \Phase1Cnt_RNO_0[6]_net_1\, N_30, N_45, 
        \Phase1Cnt[5]_net_1\, N_28_i_0, N_44, 
        \Phase1Cnt[4]_net_1\, N_26_i_0, \Phase1Cnt[0]_net_1\, 
        \Phase1Cnt[1]_net_1\, N_21, N_52, N_19, N_17, 
        \DelayCnt[0]_net_1\, \DelayCnt[1]_net_1\, 
        \PrState_ns_0_0_a2_1_3[2]\, \PrState_ns_0_0_a2_0[2]\, 
        N_65, N_115, \PrState_ns_0_0_0_tz[2]\, N_54, 
        \CycCnt[0]_net_1\, \PrState_ns[2]\, N_11_i, 
        \Phase1Cnt[2]_net_1\, \Phase1Cnt_RNIEKBN[2]_net_1\, N_7, 
        \Phase1Cnt[3]_net_1\, \Phase1Cnt_RNO_1[2]\, 
        \PrState_RNO_0_0[0]\, N_55, N_53, \Phase1Cnt[10]_net_1\, 
        N_51, \Phase1Cnt[9]_net_1\, N_49, \Phase1Cnt[6]_net_1\, 
        Phase1Cnt_n11, \Phase1Cnt[11]_net_1\, Phase1Cnt_n10, 
        Phase1Cnt_n9, N_23, N_14_i_0, \PrState_ns[3]\, N_6, 
        Phase1Cnt_n0, DelayCnt_n0, \PrState[4]_net_1\, \GND\, 
        \VCC\, GND_0, VCC_0 : std_logic;

begin 

    PrState_4 <= \PrState[4]_net_1\;
    PrState_0(4) <= \PrState_0[4]_net_1\;

    WFO : DFN1C0
      port map(D => \PrState[2]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => Adc_RdEn_inter);
    
    \PrState[2]\ : DFN1C0
      port map(D => \PrState_ns[2]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \PrState[2]_net_1\);
    
    \Phase1Cnt_RNO_0[6]\ : OA1C
      port map(A => \Phase1Cnt[5]_net_1\, B => N_45, C => 
        \Phase1Cnt[6]_net_1\, Y => \Phase1Cnt_RNO_0[6]_net_1\);
    
    \Phase1Cnt[4]\ : DFN1C0
      port map(D => N_28_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[4]_net_1\);
    
    \DelayCnt_RNO_0[4]\ : NOR2A
      port map(A => \DelayCnt[3]_net_1\, B => N_52, Y => N_55);
    
    \DelayCnt_RNIP678[1]\ : OR2B
      port map(A => \DelayCnt[1]_net_1\, B => \DelayCnt[0]_net_1\, 
        Y => N_50);
    
    \Phase1Cnt_RNO[4]\ : XA1
      port map(A => N_44, B => \Phase1Cnt[4]_net_1\, C => 
        \PrState[2]_net_1\, Y => N_28_i_0);
    
    \PrState_RNO_0[0]\ : NOR2A
      port map(A => N_54, B => \CycCnt[0]_net_1\, Y => 
        \PrState_RNO_0_0[0]\);
    
    \DelayCnt_RNIDQAC[4]\ : OR3A
      port map(A => \DelayCnt[4]_net_1\, B => \DelayCnt[2]_net_1\, 
        C => \DelayCnt[3]_net_1\, Y => 
        \PrState_ns_0_i_a2_0_0_0[1]\);
    
    \Phase1Cnt[1]\ : DFN1C0
      port map(D => N_26_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[1]_net_1\);
    
    \Phase1Cnt[11]\ : DFN1C0
      port map(D => Phase1Cnt_n11, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[11]_net_1\);
    
    \DelayCnt_RNO[1]\ : XA1
      port map(A => \DelayCnt[0]_net_1\, B => \DelayCnt[1]_net_1\, 
        C => \PrState[3]_net_1\, Y => N_17);
    
    \Phase1Cnt[5]\ : DFN1C0
      port map(D => N_30, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[5]_net_1\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \Phase1Cnt_RNO[2]\ : NOR2A
      port map(A => \PrState[2]_net_1\, B => N_11_i, Y => 
        \Phase1Cnt_RNO_1[2]\);
    
    \Phase1Cnt_RNI7MU61[4]\ : OR2B
      port map(A => \Phase1Cnt[4]_net_1\, B => N_44, Y => N_45);
    
    \Phase1Cnt_RNITDEJ2[10]\ : OR2A
      port map(A => \Phase1Cnt[10]_net_1\, B => N_51, Y => N_53);
    
    \CycCnt[0]\ : DFN1C0
      port map(D => N_6, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \CycCnt[0]_net_1\);
    
    \PrState_RNO_1[3]\ : NOR3
      port map(A => N_50, B => \PrState_ns_0_i_a2_0_0_0[1]\, C
         => \PrState_0[4]_net_1\, Y => N_64);
    
    \Phase1Cnt_RNO[1]\ : XA1
      port map(A => \Phase1Cnt[0]_net_1\, B => 
        \Phase1Cnt[1]_net_1\, C => \PrState[2]_net_1\, Y => 
        N_26_i_0);
    
    \Phase1Cnt_RNIA35V[3]\ : NOR2B
      port map(A => \Phase1Cnt[3]_net_1\, B => 
        \Phase1Cnt_RNIEKBN[2]_net_1\, Y => N_44);
    
    \Phase1Cnt_RNI5A662[8]\ : OR2B
      port map(A => \Phase1Cnt[8]_net_1\, B => N_48, Y => N_49);
    
    \PrState[1]\ : DFN1C0
      port map(D => \PrState_ns[3]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \PrState[1]_net_1\);
    
    \DelayCnt_RNO[4]\ : XA1
      port map(A => \DelayCnt[4]_net_1\, B => N_55, C => 
        \PrState[3]_net_1\, Y => N_23);
    
    \Phase1Cnt_RNO[6]\ : NOR3A
      port map(A => \PrState[2]_net_1\, B => 
        \Phase1Cnt_RNO_0[6]_net_1\, C => N_47, Y => N_32);
    
    \DelayCnt_RNI7QAC[2]\ : OR2A
      port map(A => \DelayCnt[2]_net_1\, B => N_50, Y => N_52);
    
    \Phase1Cnt_RNIEKBN[2]\ : NOR3C
      port map(A => \Phase1Cnt[0]_net_1\, B => 
        \Phase1Cnt[1]_net_1\, C => \Phase1Cnt[2]_net_1\, Y => 
        \Phase1Cnt_RNIEKBN[2]_net_1\);
    
    \PrState_RNO_0[2]\ : AOI1B
      port map(A => N_54, B => \CycCnt[0]_net_1\, C => 
        \PrState_ns_0_0_a2_1_3[2]\, Y => \PrState_ns_0_0_0_tz[2]\);
    
    \PrState_RNO[2]\ : AO1C
      port map(A => \PrState_ns_0_0_0_tz[2]\, B => RowReadOutEn, 
        C => N_65, Y => \PrState_ns[2]\);
    
    \Phase1Cnt_RNI47CU1[7]\ : NOR2B
      port map(A => \Phase1Cnt[7]_net_1\, B => N_47, Y => N_48);
    
    \CycCnt_RNO[0]\ : XA1B
      port map(A => \CycCnt[0]_net_1\, B => N_58, C => 
        \PrState[4]_net_1\, Y => N_6);
    
    \DelayCnt[2]\ : DFN1C0
      port map(D => N_19, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \DelayCnt[2]_net_1\);
    
    \PrState_RNO_0[1]\ : OR3C
      port map(A => \Phase2Cnt[0]_net_1\, B => \PrState[1]_net_1\, 
        C => RowReadOutEn_0, Y => N_68);
    
    \Phase1Cnt[0]\ : DFN1C0
      port map(D => Phase1Cnt_n0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[0]_net_1\);
    
    \Phase1Cnt_RNO[8]\ : XA1
      port map(A => N_48, B => \Phase1Cnt[8]_net_1\, C => 
        \PrState[2]_net_1\, Y => N_36);
    
    \DelayCnt[1]\ : DFN1C0
      port map(D => N_17, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \DelayCnt[1]_net_1\);
    
    \Phase1Cnt_RNIKASO2[11]\ : NOR2
      port map(A => \Phase1Cnt[11]_net_1\, B => N_53, Y => N_115);
    
    \PrState_RNO_0[3]\ : NOR2
      port map(A => \PrState[4]_net_1\, B => \PrState[3]_net_1\, 
        Y => N_63);
    
    \Phase1Cnt_RNO[10]\ : XA1A
      port map(A => \Phase1Cnt[10]_net_1\, B => N_51, C => 
        \PrState[2]_net_1\, Y => Phase1Cnt_n10);
    
    \DelayCnt[3]\ : DFN1C0
      port map(D => N_21, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \DelayCnt[3]_net_1\);
    
    \PrState_RNO[1]\ : AO1B
      port map(A => \PrState_ns_0_0_a2_0[2]\, B => N_115, C => 
        N_68, Y => \PrState_ns[3]\);
    
    \PrState[4]\ : DFN1P0
      port map(D => RowReadOutEn_i, CLK => 
        PLL_Test1_0_Sys_66M_Clk, PRE => PLL_Test1_0_SysRst_O, Q
         => \PrState[4]_net_1\);
    
    \PrState_0[4]\ : DFN1P0
      port map(D => RowReadOutEn_i, CLK => 
        PLL_Test1_0_Sys_66M_Clk, PRE => PLL_Test1_0_SysRst_O, Q
         => \PrState_0[4]_net_1\);
    
    \Phase1Cnt_RNI48IM1[6]\ : NOR3B
      port map(A => \Phase1Cnt[5]_net_1\, B => 
        \Phase1Cnt[6]_net_1\, C => N_45, Y => N_47);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \Phase1Cnt_RNO[0]\ : NOR2A
      port map(A => \PrState[2]_net_1\, B => \Phase1Cnt[0]_net_1\, 
        Y => Phase1Cnt_n0);
    
    \Phase1Cnt[10]\ : DFN1C0
      port map(D => Phase1Cnt_n10, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[10]_net_1\);
    
    \DelayCnt_RNO[2]\ : XA1A
      port map(A => \DelayCnt[2]_net_1\, B => N_50, C => 
        \PrState[3]_net_1\, Y => N_19);
    
    \DelayCnt[4]\ : DFN1C0
      port map(D => N_23, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \DelayCnt[4]_net_1\);
    
    \DelayCnt_RNO[3]\ : XA1A
      port map(A => \DelayCnt[3]_net_1\, B => N_52, C => 
        \PrState[3]_net_1\, Y => N_21);
    
    \DelayCnt[0]\ : DFN1C0
      port map(D => DelayCnt_n0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \DelayCnt[0]_net_1\);
    
    \PrState[0]\ : DFN1C0
      port map(D => N_14_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \PrState[0]_net_1\);
    
    \PrState_RNIVSG9[2]\ : NOR2B
      port map(A => RowReadOutEn_0, B => \PrState[2]_net_1\, Y
         => \PrState_ns_0_0_a2_0[2]\);
    
    \Phase1Cnt[6]\ : DFN1C0
      port map(D => N_32, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[6]_net_1\);
    
    \Phase1Cnt_RNO_0[2]\ : AX1E
      port map(A => \Phase1Cnt[0]_net_1\, B => 
        \Phase1Cnt[1]_net_1\, C => \Phase1Cnt[2]_net_1\, Y => 
        N_11_i);
    
    \Phase1Cnt_RNO[7]\ : XA1
      port map(A => N_47, B => \Phase1Cnt[7]_net_1\, C => 
        \PrState[2]_net_1\, Y => N_34);
    
    \Phase1Cnt[7]\ : DFN1C0
      port map(D => N_34, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[7]_net_1\);
    
    \Phase1Cnt_RNO[9]\ : XA1A
      port map(A => \Phase1Cnt[9]_net_1\, B => N_49, C => 
        \PrState[2]_net_1\, Y => Phase1Cnt_n9);
    
    \PrState_RNO[3]\ : NOR3A
      port map(A => RowReadOutEn_0, B => N_63, C => N_64, Y => 
        N_10);
    
    \PrState_RNIQMJF[1]\ : NOR2A
      port map(A => \PrState[1]_net_1\, B => \Phase2Cnt[0]_net_1\, 
        Y => N_54);
    
    \PrState[3]\ : DFN1C0
      port map(D => N_10, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \PrState[3]_net_1\);
    
    \Phase1Cnt_RNO[3]\ : XA1
      port map(A => \Phase1Cnt_RNIEKBN[2]_net_1\, B => 
        \Phase1Cnt[3]_net_1\, C => \PrState[2]_net_1\, Y => N_7);
    
    \Phase1Cnt[9]\ : DFN1C0
      port map(D => Phase1Cnt_n9, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[9]_net_1\);
    
    \CycCnt_RNO_1[0]\ : OR2
      port map(A => \PrState[0]_net_1\, B => \Phase2Cnt[0]_net_1\, 
        Y => \CycCnt_5_i_o2_0[0]\);
    
    \PrState_RNO_1[2]\ : OR2A
      port map(A => \PrState_ns_0_0_a2_0[2]\, B => N_115, Y => 
        N_65);
    
    \PrState_RNO[0]\ : OA1
      port map(A => \PrState_RNO_0_0[0]\, B => \PrState[0]_net_1\, 
        C => RowReadOutEn, Y => N_14_i_0);
    
    \Phase1Cnt_RNI7H0E2[9]\ : OR2A
      port map(A => \Phase1Cnt[9]_net_1\, B => N_49, Y => N_51);
    
    \Phase1Cnt[3]\ : DFN1C0
      port map(D => N_7, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[3]_net_1\);
    
    \Phase1Cnt_RNO[5]\ : XA1A
      port map(A => N_45, B => \Phase1Cnt[5]_net_1\, C => 
        \PrState[2]_net_1\, Y => N_30);
    
    \CycCnt_RNO_0[0]\ : NOR3
      port map(A => \CycCnt_5_i_o2_0[0]\, B => \PrState[3]_net_1\, 
        C => \PrState[2]_net_1\, Y => N_58);
    
    \Phase1Cnt_RNO[11]\ : XA1A
      port map(A => \Phase1Cnt[11]_net_1\, B => N_53, C => 
        \PrState[2]_net_1\, Y => Phase1Cnt_n11);
    
    \PrState_RNO_2[2]\ : OR3A
      port map(A => \PrState[3]_net_1\, B => 
        \PrState_ns_0_i_a2_0_0_0[1]\, C => N_50, Y => 
        \PrState_ns_0_0_a2_1_3[2]\);
    
    \Phase2Cnt[0]\ : DFN1C0
      port map(D => N_54, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase2Cnt[0]_net_1\);
    
    \Phase1Cnt[8]\ : DFN1C0
      port map(D => N_36, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[8]_net_1\);
    
    \Phase1Cnt[2]\ : DFN1C0
      port map(D => \Phase1Cnt_RNO_1[2]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \Phase1Cnt[2]_net_1\);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    \DelayCnt_RNO[0]\ : NOR2A
      port map(A => \PrState[3]_net_1\, B => \DelayCnt[0]_net_1\, 
        Y => DelayCnt_n0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3;
use proasic3.all;

entity WaveGenSingleZ1 is

    port( PrState_4               : in    std_logic;
          PrState_0               : in    std_logic_vector(4 to 4);
          AdcCLkEn                : out   std_logic;
          PLL_Test1_0_SysRst_O    : in    std_logic;
          PLL_Test1_0_Sys_66M_Clk : in    std_logic;
          RowReadOutEn            : in    std_logic;
          RowReadOutEn_0          : in    std_logic
        );

end WaveGenSingleZ1;

architecture DEF_ARCH of WaveGenSingleZ1 is 

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NOR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component XA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OAI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component OA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \PrState_ns_0_i_0[1]\, \PrState[3]_net_1\, 
        \PrState_ns_0_i_a2_0_2[1]\, \DelayCnt[2]_net_1\, 
        \PrState_ns_0_i_a2_0_0[1]\, \DelayCnt[0]_net_1\, 
        \DelayCnt[3]_net_1\, \DelayCnt[1]_net_1\, 
        \PrState_ns_0_0_o2_7[2]\, \PrState_ns_0_0_o2_4[2]\, 
        \Phase1Cnt[0]_net_1\, \Phase1Cnt[1]_net_1\, 
        \PrState_ns_0_0_o2_6[2]\, \PrState_ns_0_0_o2_3[2]\, 
        \Phase1Cnt[8]_net_1\, \Phase1Cnt[7]_net_1\, 
        \PrState_ns_0_0_o2_5[2]\, \PrState_ns_0_0_o2_1[2]\, 
        \Phase1Cnt[4]_net_1\, \Phase1Cnt[3]_net_1\, 
        \Phase1Cnt[9]_net_1\, \Phase1Cnt[10]_net_1\, 
        \Phase1Cnt[2]_net_1\, \Phase1Cnt[11]_net_1\, 
        \Phase1Cnt[5]_net_1\, \Phase1Cnt[6]_net_1\, 
        \CycCnt_5_i_o2_0[0]\, \PrState[0]_net_1\, 
        \Phase2Cnt[0]_net_1\, N_106, \PrState[1]_net_1\, N_8, 
        N_67, N_62, \PrState[2]_net_1\, N_34, N_47, N_32, N_46, 
        N_30, N_134, N_28, N_44, N_26, N_43, N_24, N_42, N_22_i_0, 
        N_41, N_20_i_0, N_16, N_50, N_14, 
        \PrState_ns_0_0_a2_1_2[2]\, DelayCnt_n0, 
        \PrState_ns_0_0_0[2]\, \PrState_ns_0_0_a2_0_0[2]\, N_53, 
        \CycCnt[0]_net_1\, \PrState_ns[2]\, N_145, N_78, N_76, 
        N_51, N_54, N_48, Phase1Cnt_n11, Phase1Cnt_n10, 
        Phase1Cnt_n9, N_18, N_12, \PrState_ns[3]\, N_6, 
        Phase1Cnt_n0, \GND\, \VCC\, GND_0, VCC_0 : std_logic;

begin 


    WFO : DFN1C0
      port map(D => \PrState[2]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => AdcCLkEn);
    
    \PrState[2]\ : DFN1C0
      port map(D => \PrState_ns[2]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \PrState[2]_net_1\);
    
    \Phase1Cnt_RNII46Q[3]\ : NOR3A
      port map(A => \PrState_ns_0_0_o2_1[2]\, B => 
        \Phase1Cnt[4]_net_1\, C => \Phase1Cnt[3]_net_1\, Y => 
        \PrState_ns_0_0_o2_5[2]\);
    
    \Phase1Cnt_RNO_0[6]\ : AOI1
      port map(A => \Phase1Cnt[5]_net_1\, B => N_44, C => 
        \Phase1Cnt[6]_net_1\, Y => N_134);
    
    \Phase1Cnt[4]\ : DFN1C0
      port map(D => N_26, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[4]_net_1\);
    
    \Phase1Cnt_RNO[4]\ : XA1
      port map(A => N_43, B => \Phase1Cnt[4]_net_1\, C => 
        \PrState[2]_net_1\, Y => N_26);
    
    \PrState_RNO_0[0]\ : NOR2A
      port map(A => N_53, B => \CycCnt[0]_net_1\, Y => N_78);
    
    \DelayCnt_RNO_0[3]\ : NOR2B
      port map(A => N_50, B => \DelayCnt[2]_net_1\, Y => N_54);
    
    \Phase1Cnt[1]\ : DFN1C0
      port map(D => N_20_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[1]_net_1\);
    
    \Phase1Cnt[11]\ : DFN1C0
      port map(D => Phase1Cnt_n11, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[11]_net_1\);
    
    \Phase1Cnt_RNI646Q[3]\ : NOR2A
      port map(A => \Phase1Cnt[3]_net_1\, B => N_42, Y => N_43);
    
    \DelayCnt_RNO[1]\ : XA1
      port map(A => \DelayCnt[0]_net_1\, B => \DelayCnt[1]_net_1\, 
        C => \PrState[3]_net_1\, Y => N_14);
    
    \Phase1Cnt_RNIGS932[1]\ : OR3C
      port map(A => \PrState_ns_0_0_o2_6[2]\, B => 
        \PrState_ns_0_0_o2_5[2]\, C => \PrState_ns_0_0_o2_7[2]\, 
        Y => N_67);
    
    \Phase1Cnt[5]\ : DFN1C0
      port map(D => N_28, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[5]_net_1\);
    
    \Phase1Cnt_RNIS8CK1[7]\ : NOR2B
      port map(A => \Phase1Cnt[7]_net_1\, B => N_46, Y => N_47);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \Phase1Cnt_RNO[2]\ : XA1A
      port map(A => N_41, B => \Phase1Cnt[2]_net_1\, C => 
        \PrState[2]_net_1\, Y => N_22_i_0);
    
    \CycCnt[0]\ : DFN1C0
      port map(D => N_6, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \CycCnt[0]_net_1\);
    
    \Phase1Cnt_RNIB23D[6]\ : NOR2
      port map(A => \Phase1Cnt[5]_net_1\, B => 
        \Phase1Cnt[6]_net_1\, Y => \PrState_ns_0_0_o2_1[2]\);
    
    \PrState_RNO_1[3]\ : OAI1
      port map(A => \PrState[3]_net_1\, B => PrState_0(4), C => 
        RowReadOutEn_0, Y => \PrState_ns_0_i_0[1]\);
    
    \Phase1Cnt_RNO[1]\ : XA1
      port map(A => \Phase1Cnt[0]_net_1\, B => 
        \Phase1Cnt[1]_net_1\, C => \PrState[2]_net_1\, Y => 
        N_20_i_0);
    
    \Phase1Cnt_RNI3JKJ[2]\ : OR2A
      port map(A => \Phase1Cnt[2]_net_1\, B => N_41, Y => N_42);
    
    \PrState[1]\ : DFN1C0
      port map(D => \PrState_ns[3]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \PrState[1]_net_1\);
    
    \Phase1Cnt_RNO[6]\ : NOR3A
      port map(A => \PrState[2]_net_1\, B => N_134, C => N_46, Y
         => N_30);
    
    \PrState_RNO_0[2]\ : AO1B
      port map(A => \PrState_ns_0_0_a2_1_2[2]\, B => 
        \PrState_ns_0_0_a2_0_0[2]\, C => RowReadOutEn, Y => 
        \PrState_ns_0_0_0[2]\);
    
    \Phase1Cnt_RNILNQD1[6]\ : NOR3C
      port map(A => N_44, B => \Phase1Cnt[5]_net_1\, C => 
        \Phase1Cnt[6]_net_1\, Y => N_46);
    
    \Phase1Cnt_RNI4QTQ1[8]\ : OR2B
      port map(A => \Phase1Cnt[8]_net_1\, B => N_47, Y => N_48);
    
    \PrState_RNO[2]\ : AO1B
      port map(A => N_145, B => N_67, C => \PrState_ns_0_0_0[2]\, 
        Y => \PrState_ns[2]\);
    
    \CycCnt_RNO[0]\ : XA1B
      port map(A => \CycCnt[0]_net_1\, B => N_62, C => PrState_4, 
        Y => N_6);
    
    \DelayCnt[2]\ : DFN1C0
      port map(D => N_16, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \DelayCnt[2]_net_1\);
    
    \PrState_RNO_0[1]\ : OR3C
      port map(A => \Phase2Cnt[0]_net_1\, B => \PrState[1]_net_1\, 
        C => RowReadOutEn_0, Y => N_106);
    
    \Phase1Cnt_RNIRPHK[1]\ : NOR3A
      port map(A => \PrState_ns_0_0_o2_4[2]\, B => 
        \Phase1Cnt[0]_net_1\, C => \Phase1Cnt[1]_net_1\, Y => 
        \PrState_ns_0_0_o2_7[2]\);
    
    \Phase1Cnt[0]\ : DFN1C0
      port map(D => Phase1Cnt_n0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[0]_net_1\);
    
    \Phase1Cnt_RNI3UHK[7]\ : NOR3A
      port map(A => \PrState_ns_0_0_o2_3[2]\, B => 
        \Phase1Cnt[8]_net_1\, C => \Phase1Cnt[7]_net_1\, Y => 
        \PrState_ns_0_0_o2_6[2]\);
    
    \Phase1Cnt_RNO[8]\ : XA1
      port map(A => N_47, B => \Phase1Cnt[8]_net_1\, C => 
        \PrState[2]_net_1\, Y => N_34);
    
    \DelayCnt[1]\ : DFN1C0
      port map(D => N_14, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \DelayCnt[1]_net_1\);
    
    \PrState_RNO_0[3]\ : NOR3B
      port map(A => \DelayCnt[2]_net_1\, B => 
        \PrState_ns_0_i_a2_0_0[1]\, C => \DelayCnt[0]_net_1\, Y
         => \PrState_ns_0_i_a2_0_2[1]\);
    
    \PrState_RNI6NNA[1]\ : NOR2A
      port map(A => \PrState[1]_net_1\, B => \Phase2Cnt[0]_net_1\, 
        Y => N_53);
    
    \Phase1Cnt_RNO[10]\ : XA1A
      port map(A => \Phase1Cnt[10]_net_1\, B => N_51, C => 
        \PrState[2]_net_1\, Y => Phase1Cnt_n10);
    
    \DelayCnt[3]\ : DFN1C0
      port map(D => N_18, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \DelayCnt[3]_net_1\);
    
    \PrState_RNO[1]\ : AO1C
      port map(A => N_67, B => N_145, C => N_106, Y => 
        \PrState_ns[3]\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \Phase1Cnt_RNIKRE7[11]\ : NOR2B
      port map(A => \Phase1Cnt[2]_net_1\, B => 
        \Phase1Cnt[11]_net_1\, Y => \PrState_ns_0_0_o2_3[2]\);
    
    \Phase1Cnt_RNO[0]\ : NOR2A
      port map(A => \PrState[2]_net_1\, B => \Phase1Cnt[0]_net_1\, 
        Y => Phase1Cnt_n0);
    
    \Phase1Cnt_RNIALN01[4]\ : NOR2B
      port map(A => \Phase1Cnt[4]_net_1\, B => N_43, Y => N_44);
    
    \DelayCnt_RNIIAB8[3]\ : NOR2B
      port map(A => \DelayCnt[3]_net_1\, B => \DelayCnt[1]_net_1\, 
        Y => \PrState_ns_0_i_a2_0_0[1]\);
    
    \Phase1Cnt[10]\ : DFN1C0
      port map(D => Phase1Cnt_n10, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[10]_net_1\);
    
    \DelayCnt_RNO[2]\ : XA1
      port map(A => \DelayCnt[2]_net_1\, B => N_50, C => 
        \PrState[3]_net_1\, Y => N_16);
    
    \Phase1Cnt_RNIQNE7[10]\ : NOR2
      port map(A => \Phase1Cnt[9]_net_1\, B => 
        \Phase1Cnt[10]_net_1\, Y => \PrState_ns_0_0_o2_4[2]\);
    
    \DelayCnt_RNO[3]\ : XA1
      port map(A => \DelayCnt[3]_net_1\, B => N_54, C => 
        \PrState[3]_net_1\, Y => N_18);
    
    \DelayCnt[0]\ : DFN1C0
      port map(D => DelayCnt_n0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \DelayCnt[0]_net_1\);
    
    \PrState[0]\ : DFN1C0
      port map(D => N_12, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \PrState[0]_net_1\);
    
    \Phase1Cnt[6]\ : DFN1C0
      port map(D => N_30, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[6]_net_1\);
    
    \Phase1Cnt_RNO[7]\ : XA1
      port map(A => N_46, B => \Phase1Cnt[7]_net_1\, C => 
        \PrState[2]_net_1\, Y => N_32);
    
    \Phase1Cnt[7]\ : DFN1C0
      port map(D => N_32, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[7]_net_1\);
    
    \Phase1Cnt_RNO[9]\ : XA1A
      port map(A => \Phase1Cnt[9]_net_1\, B => N_48, C => 
        \PrState[2]_net_1\, Y => Phase1Cnt_n9);
    
    \PrState_RNO[3]\ : OA1C
      port map(A => \PrState_ns_0_i_a2_0_2[1]\, B => PrState_0(4), 
        C => \PrState_ns_0_i_0[1]\, Y => N_8);
    
    \PrState[3]\ : DFN1C0
      port map(D => N_8, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \PrState[3]_net_1\);
    
    \Phase1Cnt_RNO[3]\ : XA1A
      port map(A => N_42, B => \Phase1Cnt[3]_net_1\, C => 
        \PrState[2]_net_1\, Y => N_24);
    
    \Phase1Cnt[9]\ : DFN1C0
      port map(D => Phase1Cnt_n9, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[9]_net_1\);
    
    \CycCnt_RNO_1[0]\ : OR2
      port map(A => \PrState[0]_net_1\, B => \Phase2Cnt[0]_net_1\, 
        Y => \CycCnt_5_i_o2_0[0]\);
    
    \PrState_RNO_1[2]\ : OR3C
      port map(A => \PrState_ns_0_i_a2_0_0[1]\, B => 
        \DelayCnt[2]_net_1\, C => DelayCnt_n0, Y => 
        \PrState_ns_0_0_a2_1_2[2]\);
    
    \PrState_RNIFSO9[2]\ : NOR2B
      port map(A => RowReadOutEn, B => \PrState[2]_net_1\, Y => 
        N_145);
    
    \PrState_RNO[0]\ : OA1
      port map(A => N_78, B => \PrState[0]_net_1\, C => 
        RowReadOutEn, Y => N_12);
    
    \Phase1Cnt_RNI123D[1]\ : OR2B
      port map(A => \Phase1Cnt[1]_net_1\, B => 
        \Phase1Cnt[0]_net_1\, Y => N_41);
    
    \DelayCnt_RNIKU98[0]\ : NOR2A
      port map(A => \PrState[3]_net_1\, B => \DelayCnt[0]_net_1\, 
        Y => DelayCnt_n0);
    
    \Phase1Cnt_RNO_0[11]\ : OR2A
      port map(A => \Phase1Cnt[10]_net_1\, B => N_51, Y => N_76);
    
    \Phase1Cnt[3]\ : DFN1C0
      port map(D => N_24, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[3]_net_1\);
    
    \Phase1Cnt_RNO[5]\ : XA1
      port map(A => N_44, B => \Phase1Cnt[5]_net_1\, C => 
        \PrState[2]_net_1\, Y => N_28);
    
    \CycCnt_RNO_0[0]\ : NOR3
      port map(A => \CycCnt_5_i_o2_0[0]\, B => \PrState[3]_net_1\, 
        C => \PrState[2]_net_1\, Y => N_62);
    
    \Phase1Cnt_RNO[11]\ : XA1A
      port map(A => \Phase1Cnt[11]_net_1\, B => N_76, C => 
        \PrState[2]_net_1\, Y => Phase1Cnt_n11);
    
    \PrState_RNO_2[2]\ : OR2B
      port map(A => N_53, B => \CycCnt[0]_net_1\, Y => 
        \PrState_ns_0_0_a2_0_0[2]\);
    
    \Phase2Cnt[0]\ : DFN1C0
      port map(D => N_53, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase2Cnt[0]_net_1\);
    
    \DelayCnt_RNIFUA8[1]\ : NOR2B
      port map(A => \DelayCnt[1]_net_1\, B => \DelayCnt[0]_net_1\, 
        Y => N_50);
    
    \Phase1Cnt_RNIDBF12[9]\ : OR2A
      port map(A => \Phase1Cnt[9]_net_1\, B => N_48, Y => N_51);
    
    \Phase1Cnt[8]\ : DFN1C0
      port map(D => N_34, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[8]_net_1\);
    
    \Phase1Cnt[2]\ : DFN1C0
      port map(D => N_22_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[2]_net_1\);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3;
use proasic3.all;

entity WaveGenSingleZ4 is

    port( PrState_3               : in    std_logic;
          Pre_co_c                : out   std_logic;
          PLL_Test1_0_SysRst_O    : in    std_logic;
          PLL_Test1_0_Sys_66M_Clk : in    std_logic;
          RowReadOutEn            : in    std_logic;
          RowReadOutEn_0          : in    std_logic
        );

end WaveGenSingleZ4;

architecture DEF_ARCH of WaveGenSingleZ4 is 

  component AOI1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component OR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal N_87, \PrState[1]_net_1\, \Phase2Cnt[0]_net_1\, 
        \PrState_ns_0_tz[2]\, N_77, \CycCnt[0]_net_1\, 
        \DelayCnt_RNIEUV8[0]_net_1\, \PrState_ns[2]\, N_84, N_78, 
        \Phase1Cnt[1]_net_1\, \Phase1Cnt[0]_net_1\, 
        \Phase1Cnt_4[0]\, \PrState_i[2]\, \Phase1Cnt_4[1]\, 
        \PrState[3]_net_1\, \DelayCnt[0]_net_1\, 
        \PrState_RNO_3[3]\, N_80, \PrState_ns[3]\, N_88_1, 
        \CycCnt_RNO_2[0]\, \GND\, \VCC\, GND_0, VCC_0
         : std_logic;

begin 


    \PrState_RNO[2]\ : AOI1B
      port map(A => \PrState_ns_0_tz[2]\, B => RowReadOutEn, C
         => N_84, Y => \PrState_ns[2]\);
    
    \DelayCnt[0]\ : DFN1C0
      port map(D => \DelayCnt_RNIEUV8[0]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \DelayCnt[0]_net_1\);
    
    WFO : DFN1P0
      port map(D => \PrState_i[2]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, PRE => PLL_Test1_0_SysRst_O, Q
         => Pre_co_c);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    \PrState[3]\ : DFN1C0
      port map(D => \PrState_RNO_3[3]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \PrState[3]_net_1\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \PrState[1]\ : DFN1C0
      port map(D => \PrState_ns[3]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \PrState[1]_net_1\);
    
    \PrState_RNO_0[1]\ : OR3C
      port map(A => \PrState[1]_net_1\, B => \Phase2Cnt[0]_net_1\, 
        C => RowReadOutEn_0, Y => N_87);
    
    \CycCnt[0]\ : DFN1C0
      port map(D => \CycCnt_RNO_2[0]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \CycCnt[0]_net_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \PrState_RNO[1]\ : AO1C
      port map(A => N_78, B => N_88_1, C => N_87, Y => 
        \PrState_ns[3]\);
    
    \PrState_RNIE5IB[2]\ : NOR2A
      port map(A => RowReadOutEn, B => \PrState_i[2]\, Y => 
        N_88_1);
    
    \Phase1Cnt[1]\ : DFN1C0
      port map(D => \Phase1Cnt_4[1]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \Phase1Cnt[1]_net_1\);
    
    \PrState_RNO[3]\ : OA1
      port map(A => N_80, B => PrState_3, C => RowReadOutEn, Y
         => \PrState_RNO_3[3]\);
    
    \Phase1Cnt_RNO[0]\ : NOR2
      port map(A => \PrState_i[2]\, B => \Phase1Cnt[0]_net_1\, Y
         => \Phase1Cnt_4[0]\);
    
    \CycCnt_RNO[0]\ : XA1B
      port map(A => \CycCnt[0]_net_1\, B => N_77, C => PrState_3, 
        Y => \CycCnt_RNO_2[0]\);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    \Phase1Cnt_RNO[1]\ : XA1B
      port map(A => \Phase1Cnt[0]_net_1\, B => 
        \Phase1Cnt[1]_net_1\, C => \PrState_i[2]\, Y => 
        \Phase1Cnt_4[1]\);
    
    \DelayCnt_RNIEUV8[0]\ : NOR2A
      port map(A => \PrState[3]_net_1\, B => \DelayCnt[0]_net_1\, 
        Y => \DelayCnt_RNIEUV8[0]_net_1\);
    
    \PrState_RNO_1[2]\ : OR2B
      port map(A => N_88_1, B => N_78, Y => N_84);
    
    \Phase2Cnt_RNIQDJ8[0]\ : NOR2A
      port map(A => \PrState[1]_net_1\, B => \Phase2Cnt[0]_net_1\, 
        Y => N_77);
    
    \Phase1Cnt[0]\ : DFN1C0
      port map(D => \Phase1Cnt_4[0]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \Phase1Cnt[0]_net_1\);
    
    \Phase2Cnt[0]\ : DFN1C0
      port map(D => N_77, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase2Cnt[0]_net_1\);
    
    \Phase1Cnt_RNIVIB5[1]\ : OR2B
      port map(A => \Phase1Cnt[1]_net_1\, B => 
        \Phase1Cnt[0]_net_1\, Y => N_78);
    
    \PrState_RNO_0[2]\ : AO1
      port map(A => N_77, B => \CycCnt[0]_net_1\, C => 
        \DelayCnt_RNIEUV8[0]_net_1\, Y => \PrState_ns_0_tz[2]\);
    
    \PrState_RNO_0[3]\ : NOR2B
      port map(A => \PrState[3]_net_1\, B => \DelayCnt[0]_net_1\, 
        Y => N_80);
    
    \PrState[2]\ : DFN1P0
      port map(D => \PrState_ns[2]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, PRE => PLL_Test1_0_SysRst_O, Q
         => \PrState_i[2]\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3;
use proasic3.all;

entity WaveGenSingleZ2 is

    port( PrState_3               : in    std_logic;
          PrState_0               : in    std_logic_vector(4 to 4);
          Sync_X_c                : out   std_logic;
          PLL_Test1_0_SysRst_O    : in    std_logic;
          PLL_Test1_0_Sys_66M_Clk : in    std_logic;
          RowReadOutEn_0          : in    std_logic
        );

end WaveGenSingleZ2;

architecture DEF_ARCH of WaveGenSingleZ2 is 

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component OAI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component OA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \PrState_ns_i_0[1]\, \PrState[3]_net_1\, 
        \PrState_ns_tz_0[2]\, N_104, \CycCnt[0]_net_1\, 
        \Phase1Cnt_RNIQDB2[0]_net_1\, \PrState_ns_i_a3_0_2[1]\, 
        \DelayCnt[2]_net_1\, \PrState_ns_i_a3_0_0[1]\, 
        \DelayCnt[0]_net_1\, \DelayCnt[3]_net_1\, 
        \DelayCnt[1]_net_1\, \PrState_RNO_5[3]\, 
        \PrState_RNO_1[1]_net_1\, N_119, N_120, 
        \DelayCnt_RNO[2]_net_1\, N_105, \DelayCnt_RNO[1]_net_1\, 
        \PrState_ns_a3_1_2[2]\, DelayCnt_n0, \PrState_ns[2]\, 
        N_106, \PrState[1]_net_1\, \Phase2Cnt[0]_net_1\, 
        \CycCnt_RNO_4[0]\, \DelayCnt_RNO[3]_net_1\, 
        \PrState[2]_net_1\, \Phase1Cnt[0]_net_1\, \GND\, \VCC\, 
        GND_0, VCC_0 : std_logic;

begin 


    WFO : DFN1C0
      port map(D => \PrState[2]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => Sync_X_c);
    
    \PrState[2]\ : DFN1C0
      port map(D => \PrState_ns[2]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \PrState[2]_net_1\);
    
    \Phase1Cnt_RNIQDB2[0]\ : NOR2A
      port map(A => \PrState[2]_net_1\, B => \Phase1Cnt[0]_net_1\, 
        Y => \Phase1Cnt_RNIQDB2[0]_net_1\);
    
    \DelayCnt_RNO_0[3]\ : NOR2B
      port map(A => N_105, B => \DelayCnt[2]_net_1\, Y => N_106);
    
    \DelayCnt_RNO[1]\ : XA1
      port map(A => \DelayCnt[0]_net_1\, B => \DelayCnt[1]_net_1\, 
        C => \PrState[3]_net_1\, Y => \DelayCnt_RNO[1]_net_1\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \CycCnt[0]\ : DFN1C0
      port map(D => \CycCnt_RNO_4[0]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \CycCnt[0]_net_1\);
    
    \PrState_RNO_1[3]\ : OAI1
      port map(A => PrState_0(4), B => \PrState[3]_net_1\, C => 
        RowReadOutEn_0, Y => \PrState_ns_i_0[1]\);
    
    \PrState[1]\ : DFN1C0
      port map(D => \PrState_RNO_1[1]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \PrState[1]_net_1\);
    
    \PrState_RNO_0[2]\ : NOR3C
      port map(A => \PrState_ns_i_a3_0_0[1]\, B => 
        \DelayCnt[2]_net_1\, C => DelayCnt_n0, Y => 
        \PrState_ns_a3_1_2[2]\);
    
    \PrState_RNO[2]\ : OA1
      port map(A => \PrState_ns_a3_1_2[2]\, B => 
        \PrState_ns_tz_0[2]\, C => RowReadOutEn_0, Y => 
        \PrState_ns[2]\);
    
    \CycCnt_RNO[0]\ : XA1B
      port map(A => \CycCnt[0]_net_1\, B => N_104, C => PrState_3, 
        Y => \CycCnt_RNO_4[0]\);
    
    \DelayCnt[2]\ : DFN1C0
      port map(D => \DelayCnt_RNO[2]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \DelayCnt[2]_net_1\);
    
    \PrState_RNO_0[1]\ : AOI1
      port map(A => \PrState[1]_net_1\, B => \Phase2Cnt[0]_net_1\, 
        C => \PrState[2]_net_1\, Y => N_119);
    
    \Phase1Cnt[0]\ : DFN1C0
      port map(D => \Phase1Cnt_RNIQDB2[0]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \Phase1Cnt[0]_net_1\);
    
    \DelayCnt[1]\ : DFN1C0
      port map(D => \DelayCnt_RNO[1]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \DelayCnt[1]_net_1\);
    
    \PrState_RNO_0[3]\ : NOR3B
      port map(A => \DelayCnt[2]_net_1\, B => 
        \PrState_ns_i_a3_0_0[1]\, C => \DelayCnt[0]_net_1\, Y => 
        \PrState_ns_i_a3_0_2[1]\);
    
    \DelayCnt[3]\ : DFN1C0
      port map(D => \DelayCnt_RNO[3]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \DelayCnt[3]_net_1\);
    
    \PrState_RNO[1]\ : NOR3A
      port map(A => RowReadOutEn_0, B => N_119, C => N_120, Y => 
        \PrState_RNO_1[1]_net_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \DelayCnt_RNIT1IC[1]\ : NOR2B
      port map(A => \DelayCnt[1]_net_1\, B => \DelayCnt[0]_net_1\, 
        Y => N_105);
    
    \Phase2Cnt_RNIQ9B2[0]\ : NOR2A
      port map(A => \PrState[1]_net_1\, B => \Phase2Cnt[0]_net_1\, 
        Y => N_104);
    
    \DelayCnt_RNO[2]\ : XA1
      port map(A => \DelayCnt[2]_net_1\, B => N_105, C => 
        \PrState[3]_net_1\, Y => \DelayCnt_RNO[2]_net_1\);
    
    \DelayCnt_RNO[3]\ : XA1
      port map(A => \DelayCnt[3]_net_1\, B => N_106, C => 
        \PrState[3]_net_1\, Y => \DelayCnt_RNO[3]_net_1\);
    
    \DelayCnt[0]\ : DFN1C0
      port map(D => DelayCnt_n0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \DelayCnt[0]_net_1\);
    
    \DelayCnt_RNIEAL6[0]\ : NOR2A
      port map(A => \PrState[3]_net_1\, B => \DelayCnt[0]_net_1\, 
        Y => DelayCnt_n0);
    
    \PrState_RNO[3]\ : OA1C
      port map(A => \PrState_ns_i_a3_0_2[1]\, B => PrState_0(4), 
        C => \PrState_ns_i_0[1]\, Y => \PrState_RNO_5[3]\);
    
    \PrState[3]\ : DFN1C0
      port map(D => \PrState_RNO_5[3]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \PrState[3]_net_1\);
    
    \PrState_RNO_1[2]\ : AO1
      port map(A => N_104, B => \CycCnt[0]_net_1\, C => 
        \Phase1Cnt_RNIQDB2[0]_net_1\, Y => \PrState_ns_tz_0[2]\);
    
    \DelayCnt_RNI02IC[3]\ : NOR2B
      port map(A => \DelayCnt[3]_net_1\, B => \DelayCnt[1]_net_1\, 
        Y => \PrState_ns_i_a3_0_0[1]\);
    
    \PrState_RNO_1[1]\ : NOR2
      port map(A => \PrState[1]_net_1\, B => \Phase1Cnt[0]_net_1\, 
        Y => N_120);
    
    \Phase2Cnt[0]\ : DFN1C0
      port map(D => N_104, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \Phase2Cnt[0]_net_1\);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3;
use proasic3.all;

entity adcen_dly is

    port( adcen_dly_VCC     : in    std_logic;
          adcen_dly_GND     : in    std_logic;
          Adc_RdEn_inter    : in    std_logic;
          ImageOrQl         : in    std_logic;
          CMOS_DrvX_0_AdcEn : out   std_logic
        );

end adcen_dly;

architecture DEF_ARCH of adcen_dly is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component CLKDLY
    port( CLK    : in    std_logic := 'U';
          GL     : out   std_logic;
          DLYGL0 : in    std_logic := 'U';
          DLYGL1 : in    std_logic := 'U';
          DLYGL2 : in    std_logic := 'U';
          DLYGL3 : in    std_logic := 'U';
          DLYGL4 : in    std_logic := 'U'
        );
  end component;

    signal AdcRdEn_DLY, \GND\, \VCC\, GND_0, VCC_0 : std_logic;

begin 


    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    Inst1_RNI18DB : OR2A
      port map(A => AdcRdEn_DLY, B => ImageOrQl, Y => 
        CMOS_DrvX_0_AdcEn);
    
    Inst1 : CLKDLY
      port map(CLK => Adc_RdEn_inter, GL => AdcRdEn_DLY, DLYGL0
         => adcen_dly_GND, DLYGL1 => adcen_dly_GND, DLYGL2 => 
        adcen_dly_GND, DLYGL3 => adcen_dly_VCC, DLYGL4 => 
        adcen_dly_GND);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3;
use proasic3.all;

entity WaveGenSingleZ5 is

    port( PrState_3               : in    std_logic;
          NoRowSel_c              : out   std_logic;
          PLL_Test1_0_SysRst_O    : in    std_logic;
          PLL_Test1_0_Sys_66M_Clk : in    std_logic;
          RowReadOutEn            : in    std_logic;
          RowReadOutEn_0          : in    std_logic
        );

end WaveGenSingleZ5;

architecture DEF_ARCH of WaveGenSingleZ5 is 

  component AO1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component OR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal N_86, \PrState[1]_net_1\, \Phase2Cnt[0]_net_1\, 
        \PrState_ns_0_tz[2]\, N_76, \CycCnt[0]_net_1\, 
        \DelayCnt_RNIAL36[0]_net_1\, \PrState_ns[2]\, N_83, N_77, 
        \Phase1Cnt[1]_net_1\, \Phase1Cnt[0]_net_1\, 
        \Phase1Cnt_4[0]\, \PrState[2]_net_1\, \Phase1Cnt_4[1]\, 
        \PrState[3]_net_1\, \DelayCnt[0]_net_1\, 
        \PrState_RNO_2[3]\, N_79, \PrState_ns[3]\, N_87_1, 
        \CycCnt_RNO_1[0]\, \GND\, \VCC\, GND_0, VCC_0
         : std_logic;

begin 


    \PrState_RNO[2]\ : AO1B
      port map(A => \PrState_ns_0_tz[2]\, B => RowReadOutEn, C
         => N_83, Y => \PrState_ns[2]\);
    
    \DelayCnt[0]\ : DFN1C0
      port map(D => \DelayCnt_RNIAL36[0]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \DelayCnt[0]_net_1\);
    
    \PrState_RNINMM8[2]\ : NOR2B
      port map(A => \PrState[2]_net_1\, B => RowReadOutEn, Y => 
        N_87_1);
    
    \Phase1Cnt_RNI5MT4[1]\ : OR2B
      port map(A => \Phase1Cnt[1]_net_1\, B => 
        \Phase1Cnt[0]_net_1\, Y => N_77);
    
    WFO : DFN1C0
      port map(D => \PrState[2]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => NoRowSel_c);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    \PrState[3]\ : DFN1C0
      port map(D => \PrState_RNO_2[3]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \PrState[3]_net_1\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \PrState[1]\ : DFN1C0
      port map(D => \PrState_ns[3]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \PrState[1]_net_1\);
    
    \PrState_RNO_0[1]\ : OR3C
      port map(A => \PrState[1]_net_1\, B => \Phase2Cnt[0]_net_1\, 
        C => RowReadOutEn_0, Y => N_86);
    
    \CycCnt[0]\ : DFN1C0
      port map(D => \CycCnt_RNO_1[0]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \CycCnt[0]_net_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \PrState_RNO[1]\ : AO1C
      port map(A => N_77, B => N_87_1, C => N_86, Y => 
        \PrState_ns[3]\);
    
    \Phase1Cnt[1]\ : DFN1C0
      port map(D => \Phase1Cnt_4[1]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \Phase1Cnt[1]_net_1\);
    
    \PrState_RNO[3]\ : OA1
      port map(A => N_79, B => PrState_3, C => RowReadOutEn, Y
         => \PrState_RNO_2[3]\);
    
    \Phase1Cnt_RNO[0]\ : NOR2A
      port map(A => \PrState[2]_net_1\, B => \Phase1Cnt[0]_net_1\, 
        Y => \Phase1Cnt_4[0]\);
    
    \CycCnt_RNO[0]\ : XA1B
      port map(A => \CycCnt[0]_net_1\, B => N_76, C => PrState_3, 
        Y => \CycCnt_RNO_1[0]\);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    \Phase1Cnt_RNO[1]\ : XA1
      port map(A => \Phase1Cnt[0]_net_1\, B => 
        \Phase1Cnt[1]_net_1\, C => \PrState[2]_net_1\, Y => 
        \Phase1Cnt_4[1]\);
    
    \PrState_RNO_1[2]\ : OR2B
      port map(A => N_87_1, B => N_77, Y => N_83);
    
    \Phase1Cnt[0]\ : DFN1C0
      port map(D => \Phase1Cnt_4[0]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \Phase1Cnt[0]_net_1\);
    
    \Phase2Cnt_RNIM0H5[0]\ : NOR2A
      port map(A => \PrState[1]_net_1\, B => \Phase2Cnt[0]_net_1\, 
        Y => N_76);
    
    \Phase2Cnt[0]\ : DFN1C0
      port map(D => N_76, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase2Cnt[0]_net_1\);
    
    \PrState_RNO_0[2]\ : AO1
      port map(A => N_76, B => \CycCnt[0]_net_1\, C => 
        \DelayCnt_RNIAL36[0]_net_1\, Y => \PrState_ns_0_tz[2]\);
    
    \PrState_RNO_0[3]\ : NOR2B
      port map(A => \PrState[3]_net_1\, B => \DelayCnt[0]_net_1\, 
        Y => N_79);
    
    \PrState[2]\ : DFN1C0
      port map(D => \PrState_ns[2]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \PrState[2]_net_1\);
    
    \DelayCnt_RNIAL36[0]\ : NOR2A
      port map(A => \PrState[3]_net_1\, B => \DelayCnt[0]_net_1\, 
        Y => \DelayCnt_RNIAL36[0]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3;
use proasic3.all;

entity WaveGenSinglewithCycNumSel is

    port( PrState_4               : in    std_logic;
          PrState_0               : in    std_logic_vector(4 to 4);
          Clock_X_c               : out   std_logic;
          LineReadOutOk_i         : out   std_logic;
          PLL_Test1_0_SysRst_O    : in    std_logic;
          PLL_Test1_0_Sys_66M_Clk : in    std_logic;
          RowReadOutEn            : in    std_logic;
          RowReadOutEn_0          : in    std_logic
        );

end WaveGenSinglewithCycNumSel;

architecture DEF_ARCH of WaveGenSinglewithCycNumSel is 

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component XA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1D
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component XA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component INV
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AOI1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \PrState_i[0]\, \PrState[0]_net_1\, 
        \PrState_ns_0_0_a2_1_0[2]\, \PrState[3]_net_1\, 
        CycCntlde_0_a2_1, \PrState[2]_net_1\, CycCntlde_0_a2_0, 
        \Phase2Cnt[0]_net_1\, N_12, \CycCnt[0]_net_1\, 
        \CycCnt[1]_net_1\, N_14, \CycCnt[2]_net_1\, N_151, N_16, 
        \CycCnt[3]_net_1\, N_38, N_18, \CycCnt[4]_net_1\, N_39, 
        N_20, \CycCnt[5]_net_1\, N_41, N_22, N_60, N_163, 
        N_24_i_0, \CycCnt[7]_net_1\, N_26_i_0, N_91, N_62, 
        \PrState_RNO_1[2]_net_1\, \Phase1Cnt[0]_net_1\, 
        \PrState_RNO_0_0[2]\, \DelayCnt[3]_net_1\, N_64, 
        \PrState_ns[2]\, \PrState_RNO_2[2]_net_1\, N_32, 
        \DelayCnt[2]_net_1\, N_63, N_30, \DelayCnt[0]_net_1\, 
        \DelayCnt[1]_net_1\, \PrState_ns_0_0_a2_0[2]\, N_118_1, 
        N_65, \PrState_ns[3]\, NxState_0_sqmuxa, 
        \PrState_ns_0_0_a2_0_0[3]\, \PrState[1]_net_1\, CycCnt_n0, 
        \CycCnt[6]_net_1\, \CycCnt[8]_net_1\, CycCnt_n9, 
        \CycCnt[9]_net_1\, N_66, N_34, \PrState_ns[4]\, 
        \PrState_RNO_0_1[0]\, N_6, CycCnte, DelayCnt_n0, \GND\, 
        \VCC\, GND_0, VCC_0 : std_logic;

begin 


    WFO : DFN1C0
      port map(D => \PrState[2]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => Clock_X_c);
    
    \CycCnt_RNIAPAK1[6]\ : OR3C
      port map(A => \CycCnt[5]_net_1\, B => N_41, C => 
        \CycCnt[6]_net_1\, Y => N_60);
    
    \PrState[2]\ : DFN1C0
      port map(D => \PrState_ns[2]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \PrState[2]_net_1\);
    
    \PrState_RNO_3[2]\ : NOR2B
      port map(A => \PrState[3]_net_1\, B => RowReadOutEn_0, Y
         => \PrState_ns_0_0_a2_1_0[2]\);
    
    \Phase2Cnt_RNIT4E8[0]\ : OR2
      port map(A => \Phase2Cnt[0]_net_1\, B => \PrState[0]_net_1\, 
        Y => CycCntlde_0_a2_0);
    
    \CycCnt_RNO_0[6]\ : AOI1
      port map(A => N_41, B => \CycCnt[5]_net_1\, C => 
        \CycCnt[6]_net_1\, Y => N_163);
    
    \CycCnt[9]\ : DFN1E1C0
      port map(D => CycCnt_n9, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[9]_net_1\);
    
    \CycCnt_RNO[7]\ : XA1C
      port map(A => \CycCnt[7]_net_1\, B => N_60, C => 
        PrState_0(4), Y => N_24_i_0);
    
    \PrState_RNO_0[0]\ : OR2B
      port map(A => \PrState[0]_net_1\, B => RowReadOutEn, Y => 
        \PrState_RNO_0_1[0]\);
    
    \DelayCnt_RNO[1]\ : XA1
      port map(A => \DelayCnt[0]_net_1\, B => \DelayCnt[1]_net_1\, 
        C => \PrState[3]_net_1\, Y => N_30);
    
    \Phase2Cnt_RNIH76R[0]\ : AO1D
      port map(A => CycCntlde_0_a2_1, B => CycCntlde_0_a2_0, C
         => PrState_4, Y => CycCnte);
    
    \CycCnt[8]\ : DFN1E1C0
      port map(D => N_26_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[8]_net_1\);
    
    \CycCnt[5]\ : DFN1E1C0
      port map(D => N_20, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[5]_net_1\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \CycCnt_RNO[4]\ : XA1B
      port map(A => \CycCnt[4]_net_1\, B => N_39, C => 
        PrState_0(4), Y => N_18);
    
    \CycCnt[0]\ : DFN1E1C0
      port map(D => CycCnt_n0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[0]_net_1\);
    
    \CycCnt_RNO[9]\ : XA1C
      port map(A => \CycCnt[9]_net_1\, B => N_62, C => PrState_4, 
        Y => CycCnt_n9);
    
    \PrState[1]\ : DFN1C0
      port map(D => \PrState_ns[3]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \PrState[1]_net_1\);
    
    \CycCnt_RNIC0DM[2]\ : NOR2B
      port map(A => N_151, B => \CycCnt[2]_net_1\, Y => N_38);
    
    \CycCnt_RNO[6]\ : NOR3A
      port map(A => N_60, B => N_163, C => PrState_0(4), Y => 
        N_22);
    
    \CycCnt_RNO_0[8]\ : AO1A
      port map(A => N_60, B => \CycCnt[7]_net_1\, C => 
        \CycCnt[8]_net_1\, Y => N_91);
    
    WaveRdy_RNO : INV
      port map(A => \PrState[0]_net_1\, Y => \PrState_i[0]\);
    
    \PrState_RNO_0[2]\ : OR3C
      port map(A => \DelayCnt[3]_net_1\, B => N_64, C => 
        \PrState_ns_0_0_a2_1_0[2]\, Y => \PrState_RNO_0_0[2]\);
    
    \CycCnt[2]\ : DFN1E1C0
      port map(D => N_14, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[2]_net_1\);
    
    \CycCnt_RNO[3]\ : XA1B
      port map(A => \CycCnt[3]_net_1\, B => N_38, C => 
        PrState_0(4), Y => N_16);
    
    \CycCnt_RNO[2]\ : XA1B
      port map(A => \CycCnt[2]_net_1\, B => N_151, C => 
        PrState_0(4), Y => N_14);
    
    \PrState_RNO[2]\ : OR3C
      port map(A => \PrState_RNO_0_0[2]\, B => 
        \PrState_RNO_1[2]_net_1\, C => \PrState_RNO_2[2]_net_1\, 
        Y => \PrState_ns[2]\);
    
    \CycCnt_RNO[0]\ : NOR2
      port map(A => PrState_0(4), B => \CycCnt[0]_net_1\, Y => 
        CycCnt_n0);
    
    \DelayCnt[2]\ : DFN1C0
      port map(D => N_32, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \DelayCnt[2]_net_1\);
    
    \DelayCnt_RNI7UM4[1]\ : NOR2B
      port map(A => \DelayCnt[1]_net_1\, B => \DelayCnt[0]_net_1\, 
        Y => N_63);
    
    \CycCnt[6]\ : DFN1E1C0
      port map(D => N_22, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[6]_net_1\);
    
    \PrState_RNO_0[1]\ : NOR2B
      port map(A => \PrState[1]_net_1\, B => \Phase2Cnt[0]_net_1\, 
        Y => \PrState_ns_0_0_a2_0_0[3]\);
    
    \Phase1Cnt[0]\ : DFN1C0
      port map(D => NxState_0_sqmuxa, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \Phase1Cnt[0]_net_1\);
    
    \DelayCnt[1]\ : DFN1C0
      port map(D => N_30, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \DelayCnt[1]_net_1\);
    
    \CycCnt[3]\ : DFN1E1C0
      port map(D => N_16, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[3]_net_1\);
    
    \PrState_RNIU4E8[1]\ : NOR2A
      port map(A => \PrState[1]_net_1\, B => \Phase2Cnt[0]_net_1\, 
        Y => N_118_1);
    
    \DelayCnt[3]\ : DFN1C0
      port map(D => N_34, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \DelayCnt[3]_net_1\);
    
    \PrState_RNO[1]\ : OA1
      port map(A => NxState_0_sqmuxa, B => 
        \PrState_ns_0_0_a2_0_0[3]\, C => RowReadOutEn, Y => 
        \PrState_ns[3]\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \CycCnt_RNO[1]\ : XA1B
      port map(A => \CycCnt[0]_net_1\, B => \CycCnt[1]_net_1\, C
         => PrState_0(4), Y => N_12);
    
    \CycCnt[1]\ : DFN1E1C0
      port map(D => N_12, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[1]_net_1\);
    
    \DelayCnt_RNO[2]\ : XA1
      port map(A => \DelayCnt[2]_net_1\, B => N_63, C => 
        \PrState[3]_net_1\, Y => N_32);
    
    \CycCnt_RNII8ST[3]\ : NOR2B
      port map(A => N_38, B => \CycCnt[3]_net_1\, Y => N_39);
    
    \DelayCnt_RNO[3]\ : OA1
      port map(A => \DelayCnt[3]_net_1\, B => N_64, C => N_66, Y
         => N_34);
    
    \CycCnt_RNI7STE[1]\ : NOR2B
      port map(A => \CycCnt[1]_net_1\, B => \CycCnt[0]_net_1\, Y
         => N_151);
    
    \PrState_RNIS94A[1]\ : NOR2B
      port map(A => N_118_1, B => RowReadOutEn_0, Y => 
        \PrState_ns_0_0_a2_0[2]\);
    
    \DelayCnt[0]\ : DFN1C0
      port map(D => DelayCnt_n0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \DelayCnt[0]_net_1\);
    
    \PrState[0]\ : DFN1C0
      port map(D => \PrState_ns[4]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \PrState[0]_net_1\);
    
    \DelayCnt_RNICJ27[2]\ : NOR2B
      port map(A => N_63, B => \DelayCnt[2]_net_1\, Y => N_64);
    
    \CycCnt[4]\ : DFN1E1C0
      port map(D => N_18, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[4]_net_1\);
    
    \PrState_RNO[3]\ : OA1
      port map(A => N_66, B => PrState_4, C => RowReadOutEn, Y
         => N_6);
    
    WaveRdy : DFN1P0
      port map(D => \PrState_i[0]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, PRE => PLL_Test1_0_SysRst_O, Q
         => LineReadOutOk_i);
    
    \CycCnt[7]\ : DFN1E1C0
      port map(D => N_24_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[7]_net_1\);
    
    \PrState_RNIH2TA[2]\ : OR2
      port map(A => \PrState[3]_net_1\, B => \PrState[2]_net_1\, 
        Y => CycCntlde_0_a2_1);
    
    \PrState[3]\ : DFN1C0
      port map(D => N_6, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \PrState[3]_net_1\);
    
    \DelayCnt_RNIRTSE[3]\ : AOI1B
      port map(A => N_64, B => \DelayCnt[3]_net_1\, C => 
        \PrState[3]_net_1\, Y => N_66);
    
    \PrState_RNO_1[2]\ : OR3C
      port map(A => \PrState[2]_net_1\, B => \Phase1Cnt[0]_net_1\, 
        C => RowReadOutEn_0, Y => \PrState_RNO_1[2]_net_1\);
    
    \PrState_RNO[0]\ : AO1C
      port map(A => N_65, B => \PrState_ns_0_0_a2_0[2]\, C => 
        \PrState_RNO_0_1[0]\, Y => \PrState_ns[4]\);
    
    \Phase1Cnt_RNI4GC8[0]\ : NOR2A
      port map(A => \PrState[2]_net_1\, B => \Phase1Cnt[0]_net_1\, 
        Y => NxState_0_sqmuxa);
    
    \CycCnt_RNIPKB51[4]\ : NOR2B
      port map(A => N_39, B => \CycCnt[4]_net_1\, Y => N_41);
    
    \CycCnt_RNO[5]\ : XA1B
      port map(A => \CycCnt[5]_net_1\, B => N_41, C => 
        PrState_0(4), Y => N_20);
    
    \CycCnt_RNO[8]\ : NOR3B
      port map(A => N_91, B => N_62, C => PrState_0(4), Y => 
        N_26_i_0);
    
    \CycCnt_RNIBEQA2[9]\ : OR2A
      port map(A => \CycCnt[9]_net_1\, B => N_62, Y => N_65);
    
    \CycCnt_RNIVDA32[8]\ : OR3B
      port map(A => \CycCnt[7]_net_1\, B => \CycCnt[8]_net_1\, C
         => N_60, Y => N_62);
    
    \PrState_RNO_2[2]\ : OR2B
      port map(A => \PrState_ns_0_0_a2_0[2]\, B => N_65, Y => 
        \PrState_RNO_2[2]_net_1\);
    
    \Phase2Cnt[0]\ : DFN1C0
      port map(D => N_118_1, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \Phase2Cnt[0]_net_1\);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    \DelayCnt_RNO[0]\ : NOR2A
      port map(A => \PrState[3]_net_1\, B => \DelayCnt[0]_net_1\, 
        Y => DelayCnt_n0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3;
use proasic3.all;

entity WaveGenSingleZ7 is

    port( Sync_Y_c                : out   std_logic;
          PLL_Test1_0_SysRst_O    : in    std_logic;
          PLL_Test1_0_Sys_66M_Clk : in    std_logic;
          N_30                    : in    std_logic;
          Y_X_WaveEn              : in    std_logic
        );

end WaveGenSingleZ7;

architecture DEF_ARCH of WaveGenSingleZ7 is 

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component XA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OAI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \PrState_ns_i_0[2]\, N_109, \PrState[1]_net_1\, 
        \PrState_ns_i_a4_0[2]\, \PrState[2]_net_1\, 
        \PrState[3]_net_1\, \PrState_ns_a4_0_2[3]\, 
        \PrState_ns_a4_0_0[3]\, N_123, \PrState_ns_a4_0_1[3]\, 
        \Phase1Cnt[2]_net_1\, \Phase1Cnt[3]_net_1\, 
        \PrState_ns_i_a4_1_1[2]\, N_115, 
        \Phase2Cnt_RNI6C28[0]_net_1\, \CycCnt[0]_net_1\, N_118, 
        \Phase2Cnt[0]_net_1\, N_117, \PrState_RNO[2]_net_1\, 
        \CycCnt_RNO[0]_net_1\, \Phase1Cnt_RNO[2]_net_1\, N_105, 
        \Phase1Cnt_RNO[1]_net_1\, \DelayCnt[0]_net_1\, N_106, 
        \Phase1Cnt[1]_net_1\, \Phase1Cnt[0]_net_1\, 
        \Phase1Cnt_RNO[3]_net_1\, \PrState_ns[3]\, 
        \PrState_RNO[3]_net_1\, Phase1Cnt_n0, 
        \DelayCnt_RNO[0]_net_1\, \GND\, \VCC\, GND_0, VCC_0
         : std_logic;

begin 


    WFO : DFN1C0
      port map(D => \PrState[2]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => Sync_Y_c);
    
    \PrState[2]\ : DFN1C0
      port map(D => \PrState_RNO[2]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \PrState[2]_net_1\);
    
    \PrState_RNO_3[2]\ : NOR2
      port map(A => \PrState[1]_net_1\, B => \PrState[3]_net_1\, 
        Y => \PrState_ns_i_a4_1_1[2]\);
    
    \PrState_RNO_2[1]\ : OR3C
      port map(A => \PrState[1]_net_1\, B => \Phase2Cnt[0]_net_1\, 
        C => Y_X_WaveEn, Y => N_118);
    
    \Phase1Cnt[1]\ : DFN1C0
      port map(D => \Phase1Cnt_RNO[1]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \Phase1Cnt[1]_net_1\);
    
    \PrState_RNO_4[2]\ : OR2
      port map(A => \PrState[2]_net_1\, B => \PrState[3]_net_1\, 
        Y => \PrState_ns_i_a4_0[2]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \Phase1Cnt_RNO[2]\ : XA1
      port map(A => N_105, B => \Phase1Cnt[2]_net_1\, C => 
        \PrState[2]_net_1\, Y => \Phase1Cnt_RNO[2]_net_1\);
    
    \Phase1Cnt_RNIDQHC[3]\ : NOR2A
      port map(A => \Phase1Cnt[2]_net_1\, B => 
        \Phase1Cnt[3]_net_1\, Y => \PrState_ns_a4_0_0[3]\);
    
    \CycCnt[0]\ : DFN1C0
      port map(D => \CycCnt_RNO[0]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \CycCnt[0]_net_1\);
    
    \Phase1Cnt_RNO[1]\ : NOR3A
      port map(A => \PrState[2]_net_1\, B => N_123, C => N_105, Y
         => \Phase1Cnt_RNO[1]_net_1\);
    
    \PrState[1]\ : DFN1C0
      port map(D => \PrState_ns[3]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \PrState[1]_net_1\);
    
    \PrState_RNO_0[2]\ : OAI1
      port map(A => N_109, B => \PrState[1]_net_1\, C => 
        Y_X_WaveEn, Y => \PrState_ns_i_0[2]\);
    
    \PrState_RNO[2]\ : NOR3
      port map(A => \PrState_ns_i_0[2]\, B => N_117, C => N_115, 
        Y => \PrState_RNO[2]_net_1\);
    
    \CycCnt_RNO[0]\ : XA1B
      port map(A => \CycCnt[0]_net_1\, B => 
        \Phase2Cnt_RNI6C28[0]_net_1\, C => N_30, Y => 
        \CycCnt_RNO[0]_net_1\);
    
    \Phase1Cnt_RNI9AHC[1]\ : NOR2B
      port map(A => \Phase1Cnt[1]_net_1\, B => 
        \Phase1Cnt[0]_net_1\, Y => N_105);
    
    \PrState_RNO_0[1]\ : NOR2B
      port map(A => \PrState_ns_a4_0_0[3]\, B => N_123, Y => 
        \PrState_ns_a4_0_2[3]\);
    
    \Phase1Cnt[0]\ : DFN1C0
      port map(D => Phase1Cnt_n0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[0]_net_1\);
    
    \Phase1Cnt_RNI9AHC_0[1]\ : NOR2
      port map(A => \Phase1Cnt[1]_net_1\, B => 
        \Phase1Cnt[0]_net_1\, Y => N_123);
    
    \PrState_RNO[1]\ : AO1B
      port map(A => \PrState_ns_a4_0_2[3]\, B => 
        \PrState_ns_a4_0_1[3]\, C => N_118, Y => \PrState_ns[3]\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \Phase1Cnt_RNO[0]\ : NOR2A
      port map(A => \PrState[2]_net_1\, B => \Phase1Cnt[0]_net_1\, 
        Y => Phase1Cnt_n0);
    
    \DelayCnt_RNIQ8H9[0]\ : OR2B
      port map(A => \PrState[3]_net_1\, B => \DelayCnt[0]_net_1\, 
        Y => N_109);
    
    \DelayCnt[0]\ : DFN1C0
      port map(D => \DelayCnt_RNO[0]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \DelayCnt[0]_net_1\);
    
    \PrState_RNO[3]\ : OA1A
      port map(A => N_109, B => N_30, C => Y_X_WaveEn, Y => 
        \PrState_RNO[3]_net_1\);
    
    \Phase1Cnt_RNO_0[3]\ : NOR2B
      port map(A => \Phase1Cnt[2]_net_1\, B => N_105, Y => N_106);
    
    \PrState[3]\ : DFN1C0
      port map(D => \PrState_RNO[3]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \PrState[3]_net_1\);
    
    \Phase1Cnt_RNO[3]\ : XA1
      port map(A => N_106, B => \Phase1Cnt[3]_net_1\, C => 
        \PrState[2]_net_1\, Y => \Phase1Cnt_RNO[3]_net_1\);
    
    \PrState_RNO_1[2]\ : NOR3C
      port map(A => \PrState_ns_i_a4_1_1[2]\, B => 
        \PrState_ns_a4_0_0[3]\, C => N_123, Y => N_117);
    
    \Phase1Cnt[3]\ : DFN1C0
      port map(D => \Phase1Cnt_RNO[3]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \Phase1Cnt[3]_net_1\);
    
    \PrState_RNO_2[2]\ : AOI1
      port map(A => \Phase2Cnt_RNI6C28[0]_net_1\, B => 
        \CycCnt[0]_net_1\, C => \PrState_ns_i_a4_0[2]\, Y => 
        N_115);
    
    \PrState_RNO_1[1]\ : NOR2B
      port map(A => \PrState[2]_net_1\, B => Y_X_WaveEn, Y => 
        \PrState_ns_a4_0_1[3]\);
    
    \Phase2Cnt[0]\ : DFN1C0
      port map(D => \Phase2Cnt_RNI6C28[0]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \Phase2Cnt[0]_net_1\);
    
    \Phase2Cnt_RNI6C28[0]\ : NOR2A
      port map(A => \PrState[1]_net_1\, B => \Phase2Cnt[0]_net_1\, 
        Y => \Phase2Cnt_RNI6C28[0]_net_1\);
    
    \Phase1Cnt[2]\ : DFN1C0
      port map(D => \Phase1Cnt_RNO[2]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \Phase1Cnt[2]_net_1\);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    \DelayCnt_RNO[0]\ : NOR2A
      port map(A => \PrState[3]_net_1\, B => \DelayCnt[0]_net_1\, 
        Y => \DelayCnt_RNO[0]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3;
use proasic3.all;

entity WaveGenSingleZ3 is

    port( PrState_3               : in    std_logic;
          PrState_0               : in    std_logic_vector(4 to 4);
          Sh_co_c                 : out   std_logic;
          PLL_Test1_0_SysRst_O    : in    std_logic;
          PLL_Test1_0_Sys_66M_Clk : in    std_logic;
          RowReadOutEn            : in    std_logic;
          RowReadOutEn_0          : in    std_logic
        );

end WaveGenSingleZ3;

architecture DEF_ARCH of WaveGenSingleZ3 is 

  component INV
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component XA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OAI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \PrState_i[2]\, \PrState[2]_net_1\, 
        \PrState_ns_i_0[2]\, N_109, \PrState[1]_net_1\, 
        \PrState_ns_i_a4_0[2]\, \PrState[3]_net_1\, 
        \PrState_ns_a4_0_3_1[3]\, \Phase1Cnt[1]_net_1\, 
        \PrState_ns_i_a4_1_0[2]\, \Phase1Cnt[3]_net_1\, 
        \Phase1Cnt[2]_net_1\, \PrState_ns_i_a4_1_2[2]\, 
        \Phase1Cnt[0]_net_1\, \PrState_ns_i_a4_1_1[2]\, N_116, 
        \Phase2Cnt_RNI26E3[0]_net_1\, \CycCnt[0]_net_1\, N_118, 
        \PrState_RNO_0[2]_net_1\, \CycCnt_RNO_3[0]\, 
        \Phase1Cnt_RNO_0[2]\, N_106, \Phase1Cnt_RNO_0[1]\, 
        \PrState_ns_a4_0_3[3]\, \PrState_ns[3]\, 
        \PrState_ns_a4_0[3]\, \Phase2Cnt[0]_net_1\, 
        \DelayCnt[0]_net_1\, N_107, \Phase1Cnt_RNO_0[3]_net_1\, 
        \PrState_RNO_4[3]\, Phase1Cnt_n0, \DelayCnt_RNO_0[0]\, 
        \GND\, \VCC\, GND_0, VCC_0 : std_logic;

begin 


    WFO_RNO : INV
      port map(A => \PrState[2]_net_1\, Y => \PrState_i[2]\);
    
    WFO : DFN1P0
      port map(D => \PrState_i[2]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, PRE => PLL_Test1_0_SysRst_O, Q
         => Sh_co_c);
    
    \PrState[2]\ : DFN1C0
      port map(D => \PrState_RNO_0[2]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \PrState[2]_net_1\);
    
    \PrState_RNO_3[2]\ : NOR2
      port map(A => \Phase1Cnt[1]_net_1\, B => \PrState[1]_net_1\, 
        Y => \PrState_ns_i_a4_1_1[2]\);
    
    \PrState_RNO_2[1]\ : NOR2A
      port map(A => \PrState[2]_net_1\, B => \Phase1Cnt[1]_net_1\, 
        Y => \PrState_ns_a4_0_3_1[3]\);
    
    \Phase1Cnt[1]\ : DFN1C0
      port map(D => \Phase1Cnt_RNO_0[1]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \Phase1Cnt[1]_net_1\);
    
    \PrState_RNO_4[2]\ : NOR2A
      port map(A => \Phase1Cnt[0]_net_1\, B => \PrState[3]_net_1\, 
        Y => \PrState_ns_i_a4_1_2[2]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \Phase1Cnt_RNO[2]\ : XA1
      port map(A => N_106, B => \Phase1Cnt[2]_net_1\, C => 
        \PrState[2]_net_1\, Y => \Phase1Cnt_RNO_0[2]\);
    
    \CycCnt[0]\ : DFN1C0
      port map(D => \CycCnt_RNO_3[0]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \CycCnt[0]_net_1\);
    
    \Phase1Cnt_RNO[1]\ : XA1
      port map(A => \Phase1Cnt[0]_net_1\, B => 
        \Phase1Cnt[1]_net_1\, C => \PrState[2]_net_1\, Y => 
        \Phase1Cnt_RNO_0[1]\);
    
    \PrState[1]\ : DFN1C0
      port map(D => \PrState_ns[3]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \PrState[1]_net_1\);
    
    \PrState_RNO_0[2]\ : OAI1
      port map(A => N_109, B => \PrState[1]_net_1\, C => 
        RowReadOutEn_0, Y => \PrState_ns_i_0[2]\);
    
    \PrState_RNO[2]\ : NOR3
      port map(A => \PrState_ns_i_0[2]\, B => N_118, C => N_116, 
        Y => \PrState_RNO_0[2]_net_1\);
    
    \CycCnt_RNO[0]\ : XA1B
      port map(A => \CycCnt[0]_net_1\, B => 
        \Phase2Cnt_RNI26E3[0]_net_1\, C => PrState_0(4), Y => 
        \CycCnt_RNO_3[0]\);
    
    \PrState_RNO_0[1]\ : NOR2B
      port map(A => \PrState[1]_net_1\, B => \Phase2Cnt[0]_net_1\, 
        Y => \PrState_ns_a4_0[3]\);
    
    \Phase1Cnt[0]\ : DFN1C0
      port map(D => Phase1Cnt_n0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[0]_net_1\);
    
    \PrState_RNO[1]\ : OA1
      port map(A => \PrState_ns_a4_0[3]\, B => 
        \PrState_ns_a4_0_3[3]\, C => RowReadOutEn, Y => 
        \PrState_ns[3]\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \Phase1Cnt_RNO[0]\ : NOR2A
      port map(A => \PrState[2]_net_1\, B => \Phase1Cnt[0]_net_1\, 
        Y => Phase1Cnt_n0);
    
    \Phase1Cnt_RNI7S56[3]\ : NOR2B
      port map(A => \Phase1Cnt[3]_net_1\, B => 
        \Phase1Cnt[2]_net_1\, Y => \PrState_ns_i_a4_1_0[2]\);
    
    \DelayCnt[0]\ : DFN1C0
      port map(D => \DelayCnt_RNO_0[0]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \DelayCnt[0]_net_1\);
    
    \PrState_RNO_5[2]\ : OR2
      port map(A => \PrState[2]_net_1\, B => \PrState[3]_net_1\, 
        Y => \PrState_ns_i_a4_0[2]\);
    
    \PrState_RNO[3]\ : OA1A
      port map(A => N_109, B => PrState_3, C => RowReadOutEn, Y
         => \PrState_RNO_4[3]\);
    
    \Phase1Cnt_RNO_0[3]\ : NOR2B
      port map(A => \Phase1Cnt[2]_net_1\, B => N_106, Y => N_107);
    
    \PrState[3]\ : DFN1C0
      port map(D => \PrState_RNO_4[3]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \PrState[3]_net_1\);
    
    \Phase1Cnt_RNO[3]\ : XA1
      port map(A => N_107, B => \Phase1Cnt[3]_net_1\, C => 
        \PrState[2]_net_1\, Y => \Phase1Cnt_RNO_0[3]_net_1\);
    
    \Phase1Cnt_RNI3S56[1]\ : NOR2B
      port map(A => \Phase1Cnt[1]_net_1\, B => 
        \Phase1Cnt[0]_net_1\, Y => N_106);
    
    \DelayCnt_RNIAEI4[0]\ : OR2B
      port map(A => \PrState[3]_net_1\, B => \DelayCnt[0]_net_1\, 
        Y => N_109);
    
    \PrState_RNO_1[2]\ : NOR3C
      port map(A => \PrState_ns_i_a4_1_1[2]\, B => 
        \PrState_ns_i_a4_1_0[2]\, C => \PrState_ns_i_a4_1_2[2]\, 
        Y => N_118);
    
    \Phase1Cnt[3]\ : DFN1C0
      port map(D => \Phase1Cnt_RNO_0[3]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \Phase1Cnt[3]_net_1\);
    
    \PrState_RNO_2[2]\ : AOI1
      port map(A => \Phase2Cnt_RNI26E3[0]_net_1\, B => 
        \CycCnt[0]_net_1\, C => \PrState_ns_i_a4_0[2]\, Y => 
        N_116);
    
    \PrState_RNO_1[1]\ : NOR3C
      port map(A => \PrState_ns_i_a4_1_0[2]\, B => 
        \Phase1Cnt[0]_net_1\, C => \PrState_ns_a4_0_3_1[3]\, Y
         => \PrState_ns_a4_0_3[3]\);
    
    \Phase2Cnt[0]\ : DFN1C0
      port map(D => \Phase2Cnt_RNI26E3[0]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \Phase2Cnt[0]_net_1\);
    
    \Phase1Cnt[2]\ : DFN1C0
      port map(D => \Phase1Cnt_RNO_0[2]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \Phase1Cnt[2]_net_1\);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    \Phase2Cnt_RNI26E3[0]\ : NOR2A
      port map(A => \PrState[1]_net_1\, B => \Phase2Cnt[0]_net_1\, 
        Y => \Phase2Cnt_RNI26E3[0]_net_1\);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    \DelayCnt_RNO[0]\ : NOR2A
      port map(A => \PrState[3]_net_1\, B => \DelayCnt[0]_net_1\, 
        Y => \DelayCnt_RNO_0[0]\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3;
use proasic3.all;

entity Y_X_Addressing is

    port( Clock_X_c               : out   std_logic;
          Sync_X_c                : out   std_logic;
          Sh_co_c                 : out   std_logic;
          Pre_co_c                : out   std_logic;
          NoRowSel_c              : out   std_logic;
          Clock_Y_c               : out   std_logic;
          Sync_Y_c                : out   std_logic;
          CMOS_DrvX_0_AdcEn       : out   std_logic;
          ImageOrQl               : in    std_logic;
          DRY_c_c                 : out   std_logic;
          PLL_Test1_0_ADC_66M_Clk : in    std_logic;
          Y_X_Addressing_GND      : in    std_logic;
          Y_X_Addressing_VCC      : in    std_logic;
          Y_X_WaveEn_i            : in    std_logic;
          Y_X_WaveOk              : out   std_logic;
          Y_X_WaveEn              : in    std_logic;
          PLL_Test1_0_SysRst_O    : in    std_logic;
          PLL_Test1_0_Sys_66M_Clk : in    std_logic
        );

end Y_X_Addressing;

architecture DEF_ARCH of Y_X_Addressing is 

  component DFN1E1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component WaveGenSingleZ6
    port( PrState_3               : in    std_logic := 'U';
          Clock_Y_c               : out   std_logic;
          PLL_Test1_0_SysRst_O    : in    std_logic := 'U';
          PLL_Test1_0_Sys_66M_Clk : in    std_logic := 'U';
          RowReadOutEn            : in    std_logic := 'U';
          RowReadOutEn_0          : in    std_logic := 'U'
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component AOI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component sampleEn_dly
    port( sampleEn_dly_VCC        : in    std_logic := 'U';
          sampleEn_dly_GND        : in    std_logic := 'U';
          AdcCLkEn                : in    std_logic := 'U';
          PLL_Test1_0_ADC_66M_Clk : in    std_logic := 'U';
          DRY_c_c                 : out   std_logic
        );
  end component;

  component XA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component WaveGenSingleZ0
    port( PrState_4               : out   std_logic;
          PrState_0               : out   std_logic_vector(4 to 4);
          Adc_RdEn_inter          : out   std_logic;
          RowReadOutEn            : in    std_logic := 'U';
          RowReadOutEn_0          : in    std_logic := 'U';
          PLL_Test1_0_SysRst_O    : in    std_logic := 'U';
          RowReadOutEn_i          : in    std_logic := 'U';
          PLL_Test1_0_Sys_66M_Clk : in    std_logic := 'U'
        );
  end component;

  component WaveGenSingleZ1
    port( PrState_4               : in    std_logic := 'U';
          PrState_0               : in    std_logic_vector(4 to 4) := (others => 'U');
          AdcCLkEn                : out   std_logic;
          PLL_Test1_0_SysRst_O    : in    std_logic := 'U';
          PLL_Test1_0_Sys_66M_Clk : in    std_logic := 'U';
          RowReadOutEn            : in    std_logic := 'U';
          RowReadOutEn_0          : in    std_logic := 'U'
        );
  end component;

  component WaveGenSingleZ4
    port( PrState_3               : in    std_logic := 'U';
          Pre_co_c                : out   std_logic;
          PLL_Test1_0_SysRst_O    : in    std_logic := 'U';
          PLL_Test1_0_Sys_66M_Clk : in    std_logic := 'U';
          RowReadOutEn            : in    std_logic := 'U';
          RowReadOutEn_0          : in    std_logic := 'U'
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component WaveGenSingleZ2
    port( PrState_3               : in    std_logic := 'U';
          PrState_0               : in    std_logic_vector(4 to 4) := (others => 'U');
          Sync_X_c                : out   std_logic;
          PLL_Test1_0_SysRst_O    : in    std_logic := 'U';
          PLL_Test1_0_Sys_66M_Clk : in    std_logic := 'U';
          RowReadOutEn_0          : in    std_logic := 'U'
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component adcen_dly
    port( adcen_dly_VCC     : in    std_logic := 'U';
          adcen_dly_GND     : in    std_logic := 'U';
          Adc_RdEn_inter    : in    std_logic := 'U';
          ImageOrQl         : in    std_logic := 'U';
          CMOS_DrvX_0_AdcEn : out   std_logic
        );
  end component;

  component NOR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component WaveGenSingleZ5
    port( PrState_3               : in    std_logic := 'U';
          NoRowSel_c              : out   std_logic;
          PLL_Test1_0_SysRst_O    : in    std_logic := 'U';
          PLL_Test1_0_Sys_66M_Clk : in    std_logic := 'U';
          RowReadOutEn            : in    std_logic := 'U';
          RowReadOutEn_0          : in    std_logic := 'U'
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component INV
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component WaveGenSinglewithCycNumSel
    port( PrState_4               : in    std_logic := 'U';
          PrState_0               : in    std_logic_vector(4 to 4) := (others => 'U');
          Clock_X_c               : out   std_logic;
          LineReadOutOk_i         : out   std_logic;
          PLL_Test1_0_SysRst_O    : in    std_logic := 'U';
          PLL_Test1_0_Sys_66M_Clk : in    std_logic := 'U';
          RowReadOutEn            : in    std_logic := 'U';
          RowReadOutEn_0          : in    std_logic := 'U'
        );
  end component;

  component OR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component WaveGenSingleZ7
    port( Sync_Y_c                : out   std_logic;
          PLL_Test1_0_SysRst_O    : in    std_logic := 'U';
          PLL_Test1_0_Sys_66M_Clk : in    std_logic := 'U';
          N_30                    : in    std_logic := 'U';
          Y_X_WaveEn              : in    std_logic := 'U'
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component WaveGenSingleZ3
    port( PrState_3               : in    std_logic := 'U';
          PrState_0               : in    std_logic_vector(4 to 4) := (others => 'U');
          Sh_co_c                 : out   std_logic;
          PLL_Test1_0_SysRst_O    : in    std_logic := 'U';
          PLL_Test1_0_Sys_66M_Clk : in    std_logic := 'U';
          RowReadOutEn            : in    std_logic := 'U';
          RowReadOutEn_0          : in    std_logic := 'U'
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \RowReadOutEn_0\, \PrState[3]_net_1\, RowReadOutEn_i, 
        \PrState_ns_0_a3_0_0[4]\, N_171_1, RowCnt_n10_0_0_a3_0_0, 
        \RowCnt[9]_net_1\, N_30, \RowCnt[10]_net_1\, 
        RowCnt_n10_0_0_a3_0, \PrState_ns[3]\, LineReadOutOk_i, 
        \PrState[2]_net_1\, \PrState_RNO_6[3]\, N_166, N_167, 
        \PrState_RNO_3[2]\, N_168, N_25_i_0, N_73, N_162, 
        N_23_i_0, N_34, \RowCnt[7]_net_1\, N_21, N_71, N_19, N_31, 
        \RowCnt[5]_net_1\, N_17, N_160, \RowCnt[4]_net_1\, N_15, 
        N_29, \RowCnt[3]_net_1\, N_13, N_28, \RowCnt[2]_net_1\, 
        N_11, RowCnt_c0, \RowCnt[1]_net_1\, N_158, 
        \PrState[1]_net_1\, N_163, RowCnt_n10, \PrState_ns[4]\, 
        N_170, \PrState[0]_net_1\, \RowCnt[8]_net_1\, 
        \RowCnt[6]_net_1\, RowCnt_n9, RowCnt_n0, \RowReadOutEn\, 
        AdcCLkEn, Adc_RdEn_inter, \PrState[4]_net_1\, 
        \PrState_0[4]\, \GND\, \VCC\, GND_0, VCC_0 : std_logic;

    for all : WaveGenSingleZ6
	Use entity work.WaveGenSingleZ6(DEF_ARCH);
    for all : sampleEn_dly
	Use entity work.sampleEn_dly(DEF_ARCH);
    for all : WaveGenSingleZ0
	Use entity work.WaveGenSingleZ0(DEF_ARCH);
    for all : WaveGenSingleZ1
	Use entity work.WaveGenSingleZ1(DEF_ARCH);
    for all : WaveGenSingleZ4
	Use entity work.WaveGenSingleZ4(DEF_ARCH);
    for all : WaveGenSingleZ2
	Use entity work.WaveGenSingleZ2(DEF_ARCH);
    for all : adcen_dly
	Use entity work.adcen_dly(DEF_ARCH);
    for all : WaveGenSingleZ5
	Use entity work.WaveGenSingleZ5(DEF_ARCH);
    for all : WaveGenSinglewithCycNumSel
	Use entity work.WaveGenSinglewithCycNumSel(DEF_ARCH);
    for all : WaveGenSingleZ7
	Use entity work.WaveGenSingleZ7(DEF_ARCH);
    for all : WaveGenSingleZ3
	Use entity work.WaveGenSingleZ3(DEF_ARCH);
begin 


    \RowCnt[2]\ : DFN1E1C0
      port map(D => N_13, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => N_158, Q => \RowCnt[2]_net_1\);
    
    \RowCnt_RNIJ0FC[1]\ : NOR2B
      port map(A => \RowCnt[1]_net_1\, B => RowCnt_c0, Y => N_28);
    
    \PrState[2]\ : DFN1C0
      port map(D => \PrState_RNO_3[2]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \PrState[2]_net_1\);
    
    Wave_Clock_Y : WaveGenSingleZ6
      port map(PrState_3 => \PrState[4]_net_1\, Clock_Y_c => 
        Clock_Y_c, PLL_Test1_0_SysRst_O => PLL_Test1_0_SysRst_O, 
        PLL_Test1_0_Sys_66M_Clk => PLL_Test1_0_Sys_66M_Clk, 
        RowReadOutEn => \RowReadOutEn\, RowReadOutEn_0 => 
        \RowReadOutEn_0\);
    
    \RowCnt_RNO[10]\ : MX2
      port map(A => RowCnt_n10_0_0_a3_0_0, B => 
        RowCnt_n10_0_0_a3_0, S => N_163, Y => RowCnt_n10);
    
    \RowCnt[4]\ : DFN1E1C0
      port map(D => N_17, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => N_158, Q => \RowCnt[4]_net_1\);
    
    \RowCnt_RNIKIKB1[6]\ : OR3C
      port map(A => N_31, B => \RowCnt[5]_net_1\, C => 
        \RowCnt[6]_net_1\, Y => N_34);
    
    \RowCnt[9]\ : DFN1E1C0
      port map(D => RowCnt_n9, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => N_158, Q => 
        \RowCnt[9]_net_1\);
    
    \PrState_RNO_0[0]\ : NOR2B
      port map(A => Y_X_WaveEn, B => N_171_1, Y => 
        \PrState_ns_0_a3_0_0[4]\);
    
    RowReadOutEn : DFN1C0
      port map(D => \PrState[3]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \RowReadOutEn\);
    
    \RowCnt_RNO_1[10]\ : NOR2A
      port map(A => \RowCnt[10]_net_1\, B => N_30, Y => 
        RowCnt_n10_0_0_a3_0);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \RowCnt_RNO_0[6]\ : AOI1
      port map(A => \RowCnt[5]_net_1\, B => N_31, C => 
        \RowCnt[6]_net_1\, Y => N_71);
    
    ADCCLKDlYEn : sampleEn_dly
      port map(sampleEn_dly_VCC => Y_X_Addressing_VCC, 
        sampleEn_dly_GND => Y_X_Addressing_GND, AdcCLkEn => 
        AdcCLkEn, PLL_Test1_0_ADC_66M_Clk => 
        PLL_Test1_0_ADC_66M_Clk, DRY_c_c => DRY_c_c);
    
    \RowCnt_RNINH5V[4]\ : NOR2B
      port map(A => \RowCnt[4]_net_1\, B => N_160, Y => N_31);
    
    \RowCnt_RNO[9]\ : XA1C
      port map(A => \RowCnt[9]_net_1\, B => N_162, C => N_30, Y
         => RowCnt_n9);
    
    \PrState_RNO_1[3]\ : NOR2A
      port map(A => N_171_1, B => N_163, Y => N_167);
    
    ADC_RdENGen : WaveGenSingleZ0
      port map(PrState_4 => \PrState[4]_net_1\, PrState_0(4) => 
        \PrState_0[4]\, Adc_RdEn_inter => Adc_RdEn_inter, 
        RowReadOutEn => \RowReadOutEn\, RowReadOutEn_0 => 
        \RowReadOutEn_0\, PLL_Test1_0_SysRst_O => 
        PLL_Test1_0_SysRst_O, RowReadOutEn_i => RowReadOutEn_i, 
        PLL_Test1_0_Sys_66M_Clk => PLL_Test1_0_Sys_66M_Clk);
    
    ADC_Clock_EN : WaveGenSingleZ1
      port map(PrState_4 => \PrState[4]_net_1\, PrState_0(4) => 
        \PrState_0[4]\, AdcCLkEn => AdcCLkEn, 
        PLL_Test1_0_SysRst_O => PLL_Test1_0_SysRst_O, 
        PLL_Test1_0_Sys_66M_Clk => PLL_Test1_0_Sys_66M_Clk, 
        RowReadOutEn => \RowReadOutEn\, RowReadOutEn_0 => 
        \RowReadOutEn_0\);
    
    Wave_Pre_co : WaveGenSingleZ4
      port map(PrState_3 => \PrState[4]_net_1\, Pre_co_c => 
        Pre_co_c, PLL_Test1_0_SysRst_O => PLL_Test1_0_SysRst_O, 
        PLL_Test1_0_Sys_66M_Clk => PLL_Test1_0_Sys_66M_Clk, 
        RowReadOutEn => \RowReadOutEn\, RowReadOutEn_0 => 
        \RowReadOutEn_0\);
    
    \RowCnt_RNI74BU1[9]\ : OR2A
      port map(A => \RowCnt[9]_net_1\, B => N_162, Y => N_163);
    
    \PrState[1]\ : DFN1C0
      port map(D => \PrState_ns[3]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \PrState[1]_net_1\);
    
    \RowCnt[8]\ : DFN1E1C0
      port map(D => N_25_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => N_158, Q => 
        \RowCnt[8]_net_1\);
    
    \RowCnt[3]\ : DFN1E1C0
      port map(D => N_15, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => N_158, Q => \RowCnt[3]_net_1\);
    
    \RowCnt[10]\ : DFN1E1C0
      port map(D => RowCnt_n10, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => N_158, Q => 
        \RowCnt[10]_net_1\);
    
    Wave_Sync_X : WaveGenSingleZ2
      port map(PrState_3 => \PrState[4]_net_1\, PrState_0(4) => 
        \PrState_0[4]\, Sync_X_c => Sync_X_c, 
        PLL_Test1_0_SysRst_O => PLL_Test1_0_SysRst_O, 
        PLL_Test1_0_Sys_66M_Clk => PLL_Test1_0_Sys_66M_Clk, 
        RowReadOutEn_0 => \RowReadOutEn_0\);
    
    \PrState_RNO_0[2]\ : NOR2
      port map(A => \PrState[3]_net_1\, B => \PrState[2]_net_1\, 
        Y => N_168);
    
    \PrState_RNIBPB5[1]\ : OR2
      port map(A => \PrState[1]_net_1\, B => N_30, Y => N_158);
    
    \RowCnt_RNO_0[8]\ : AO1A
      port map(A => N_34, B => \RowCnt[7]_net_1\, C => 
        \RowCnt[8]_net_1\, Y => N_73);
    
    \RowCnt_RNO[2]\ : XA1B
      port map(A => N_28, B => \RowCnt[2]_net_1\, C => N_30, Y
         => N_13);
    
    \RowCnt_RNO[1]\ : XA1B
      port map(A => RowCnt_c0, B => \RowCnt[1]_net_1\, C => N_30, 
        Y => N_11);
    
    ADCrdDlYEn : adcen_dly
      port map(adcen_dly_VCC => Y_X_Addressing_VCC, adcen_dly_GND
         => Y_X_Addressing_GND, Adc_RdEn_inter => Adc_RdEn_inter, 
        ImageOrQl => ImageOrQl, CMOS_DrvX_0_AdcEn => 
        CMOS_DrvX_0_AdcEn);
    
    \PrState_RNO[2]\ : NOR3A
      port map(A => Y_X_WaveEn, B => N_168, C => LineReadOutOk_i, 
        Y => \PrState_RNO_3[2]\);
    
    \Y_X_WaveOk\ : DFN1C0
      port map(D => \PrState[0]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => Y_X_WaveOk);
    
    \RowCnt_RNO[4]\ : XA1B
      port map(A => N_160, B => \RowCnt[4]_net_1\, C => N_30, Y
         => N_17);
    
    \PrState_RNO_0[3]\ : AOI1
      port map(A => \PrState[3]_net_1\, B => LineReadOutOk_i, C
         => N_158, Y => N_166);
    
    Wave_NoRowSel : WaveGenSingleZ5
      port map(PrState_3 => \PrState[4]_net_1\, NoRowSel_c => 
        NoRowSel_c, PLL_Test1_0_SysRst_O => PLL_Test1_0_SysRst_O, 
        PLL_Test1_0_Sys_66M_Clk => PLL_Test1_0_Sys_66M_Clk, 
        RowReadOutEn => \RowReadOutEn\, RowReadOutEn_0 => 
        \RowReadOutEn_0\);
    
    \PrState_RNO[1]\ : NOR3C
      port map(A => LineReadOutOk_i, B => \PrState[2]_net_1\, C
         => Y_X_WaveEn, Y => \PrState_ns[3]\);
    
    \PrState[4]\ : DFN1P0
      port map(D => Y_X_WaveEn_i, CLK => PLL_Test1_0_Sys_66M_Clk, 
        PRE => PLL_Test1_0_SysRst_O, Q => N_30);
    
    GND_i : GND
      port map(Y => \GND\);
    
    RowReadOutEn_0_RNIU4M1 : INV
      port map(A => \RowReadOutEn_0\, Y => RowReadOutEn_i);
    
    \RowCnt[6]\ : DFN1E1C0
      port map(D => N_21, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => N_158, Q => \RowCnt[6]_net_1\);
    
    \RowCnt[5]\ : DFN1E1C0
      port map(D => N_19, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => N_158, Q => \RowCnt[5]_net_1\);
    
    \RowCnt_RNIA1UO[3]\ : NOR2B
      port map(A => \RowCnt[3]_net_1\, B => N_29, Y => N_160);
    
    \PrState[0]\ : DFN1C0
      port map(D => \PrState_ns[4]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \PrState[0]_net_1\);
    
    Wave_Clock_X : WaveGenSinglewithCycNumSel
      port map(PrState_4 => \PrState[4]_net_1\, PrState_0(4) => 
        \PrState_0[4]\, Clock_X_c => Clock_X_c, LineReadOutOk_i
         => LineReadOutOk_i, PLL_Test1_0_SysRst_O => 
        PLL_Test1_0_SysRst_O, PLL_Test1_0_Sys_66M_Clk => 
        PLL_Test1_0_Sys_66M_Clk, RowReadOutEn => \RowReadOutEn\, 
        RowReadOutEn_0 => \RowReadOutEn_0\);
    
    \RowCnt_RNIUGMI[2]\ : NOR2B
      port map(A => \RowCnt[2]_net_1\, B => N_28, Y => N_29);
    
    \RowCnt_RNILJ3O1[8]\ : OR3B
      port map(A => \RowCnt[7]_net_1\, B => \RowCnt[8]_net_1\, C
         => N_34, Y => N_162);
    
    \RowCnt[1]\ : DFN1E1C0
      port map(D => N_11, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => N_158, Q => \RowCnt[1]_net_1\);
    
    RowReadOutEn_0 : DFN1C0
      port map(D => \PrState[3]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \RowReadOutEn_0\);
    
    \PrState_RNIEOE4[1]\ : NOR2B
      port map(A => \RowCnt[10]_net_1\, B => \PrState[1]_net_1\, 
        Y => N_171_1);
    
    \RowCnt_RNO_0[10]\ : NOR3A
      port map(A => \RowCnt[9]_net_1\, B => N_30, C => 
        \RowCnt[10]_net_1\, Y => RowCnt_n10_0_0_a3_0_0);
    
    \PrState_RNO[3]\ : NOR3A
      port map(A => Y_X_WaveEn, B => N_166, C => N_167, Y => 
        \PrState_RNO_6[3]\);
    
    Wave_Sync_Y : WaveGenSingleZ7
      port map(Sync_Y_c => Sync_Y_c, PLL_Test1_0_SysRst_O => 
        PLL_Test1_0_SysRst_O, PLL_Test1_0_Sys_66M_Clk => 
        PLL_Test1_0_Sys_66M_Clk, N_30 => N_30, Y_X_WaveEn => 
        Y_X_WaveEn);
    
    \RowCnt[7]\ : DFN1E1C0
      port map(D => N_23_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => N_158, Q => 
        \RowCnt[7]_net_1\);
    
    \PrState[3]\ : DFN1C0
      port map(D => \PrState_RNO_6[3]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \PrState[3]_net_1\);
    
    \RowCnt_RNO[6]\ : NOR3A
      port map(A => N_34, B => N_71, C => N_30, Y => N_21);
    
    \RowCnt_RNO[8]\ : NOR3B
      port map(A => N_73, B => N_162, C => N_30, Y => N_25_i_0);
    
    \RowCnt_RNO[0]\ : NOR2
      port map(A => RowCnt_c0, B => N_30, Y => RowCnt_n0);
    
    \PrState_RNO[0]\ : AO1C
      port map(A => N_163, B => \PrState_ns_0_a3_0_0[4]\, C => 
        N_170, Y => \PrState_ns[4]\);
    
    Wave_Sh_co : WaveGenSingleZ3
      port map(PrState_3 => \PrState[4]_net_1\, PrState_0(4) => 
        \PrState_0[4]\, Sh_co_c => Sh_co_c, PLL_Test1_0_SysRst_O
         => PLL_Test1_0_SysRst_O, PLL_Test1_0_Sys_66M_Clk => 
        PLL_Test1_0_Sys_66M_Clk, RowReadOutEn => \RowReadOutEn\, 
        RowReadOutEn_0 => \RowReadOutEn_0\);
    
    \RowCnt_RNO[7]\ : XA1C
      port map(A => N_34, B => \RowCnt[7]_net_1\, C => N_30, Y
         => N_23_i_0);
    
    \RowCnt_RNO[3]\ : XA1B
      port map(A => N_29, B => \RowCnt[3]_net_1\, C => N_30, Y
         => N_15);
    
    \RowCnt[0]\ : DFN1E1C0
      port map(D => RowCnt_n0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => N_158, Q => RowCnt_c0);
    
    \RowCnt_RNO[5]\ : XA1B
      port map(A => N_31, B => \RowCnt[5]_net_1\, C => N_30, Y
         => N_19);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    \PrState_RNO_1[0]\ : OR2B
      port map(A => Y_X_WaveEn, B => \PrState[0]_net_1\, Y => 
        N_170);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3;
use proasic3.all;

entity CMOS_Ctl is

    port( CMOS_Ctl_GND             : in    std_logic;
          CMOS_DrvX_0_SDramEn      : out   std_logic;
          ImageOrQl                : out   std_logic;
          SPI_En                   : out   std_logic;
          PAT_En                   : out   std_logic;
          CMOS_DrvX_0_LVDSen       : out   std_logic;
          FrameMk_0_LVDS_ok        : in    std_logic;
          Sdram_cmd_0_SDoneFrameOk : in    std_logic;
          Y_X_WaveOk               : in    std_logic;
          PAT_Ok                   : in    std_logic;
          SPI_Ok                   : in    std_logic;
          SPI_En_i                 : out   std_logic;
          Y_X_WaveEn               : out   std_logic;
          Y_X_WaveEn_i             : out   std_logic;
          SPI_En_0                 : out   std_logic;
          CMOS_DrvX_0_SDramEn_0    : out   std_logic;
          CMOS_DrvX_0_SDramEn_1    : out   std_logic;
          CMOS_DrvX_0_SDramEn_2    : out   std_logic;
          CMOS_DrvX_0_SDramEn_3    : out   std_logic;
          CMOS_DrvX_0_SDramEn_4    : out   std_logic;
          CMOS_DrvX_0_SDramEn_5    : out   std_logic;
          CMOS_DrvX_0_LVDSen_0     : out   std_logic;
          CMOS_DrvX_0_LVDSen_1     : out   std_logic;
          CMOS_DrvX_0_LVDSen_2     : out   std_logic;
          PLL_Test1_0_SysRst_O     : in    std_logic;
          PLL_Test1_0_Sys_66M_Clk  : in    std_logic;
          CMOS_DrvX_0_LVDSen_3     : out   std_logic
        );

end CMOS_Ctl;

architecture DEF_ARCH of CMOS_Ctl is 

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component XA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E0C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component INV
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component NOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \PrState[0]_net_1\, \PrState_RNI9G29[2]_net_1\, 
        \PrState[5]_net_1\, SPI_En_0_net_1, \PrState_ns_1[3]\, 
        N_115, N_114, N_117, \PrState_ns_0_a3_0_2[7]\, 
        \PrState[1]_net_1\, \ACCcnt[5]_net_1\, \ACCcnt[4]_net_1\, 
        \PrState_ns_0_a3_0_1[7]\, \ACCcnt[2]_net_1\, 
        \ACCcnt[3]_net_1\, N_27_i_0, N_32, N_15, N_20, N_13, N_19, 
        N_128, N_18, N_127, \PrState_ns[3]\, N_21, 
        \ACCcnt[1]_net_1\, \ACCcnt[0]_net_1\, N_17, ACCcnt_n0, 
        N_124, N_112, \PrState[4]_net_1\, N_118, 
        \PrState[3]_net_1\, N_120, \PrState[2]_net_1\, 
        \Y_X_WaveEn_RNO\, \PrState[6]_net_1\, \PrState_ns[1]\, 
        \PrState[7]_net_1\, \PrState_ns[2]\, \PrState_ns[4]\, 
        \PrState_ns[5]\, \PrState_RNO[1]_net_1\, \PrState_ns[7]\, 
        Y_X_WaveEn_net_1, \GND\, \VCC\, GND_0, VCC_0 : std_logic;

begin 

    Y_X_WaveEn <= Y_X_WaveEn_net_1;
    SPI_En_0 <= SPI_En_0_net_1;

    LVDSen_2 : DFN1C0
      port map(D => \PrState[0]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => CMOS_DrvX_0_LVDSen_2);
    
    \ACCcnt_RNO[5]\ : XA1B
      port map(A => \ACCcnt[5]_net_1\, B => N_21, C => 
        \PrState[0]_net_1\, Y => N_17);
    
    \PrState[2]\ : DFN1C0
      port map(D => \PrState_ns[5]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \PrState[2]_net_1\);
    
    LVDSen_1 : DFN1C0
      port map(D => \PrState[0]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => CMOS_DrvX_0_LVDSen_1);
    
    \ACCcnt_RNIARK9[5]\ : NOR3A
      port map(A => \PrState[1]_net_1\, B => \ACCcnt[5]_net_1\, C
         => \ACCcnt[4]_net_1\, Y => \PrState_ns_0_a3_0_2[7]\);
    
    \ACCcnt_RNIVO35[1]\ : NOR2B
      port map(A => \ACCcnt[1]_net_1\, B => \ACCcnt[0]_net_1\, Y
         => N_18);
    
    \ACCcnt[1]\ : DFN1E0C0
      port map(D => N_127, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => N_124, Q => 
        \ACCcnt[1]_net_1\);
    
    SDramEn_5 : DFN1C0
      port map(D => \PrState_RNI9G29[2]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => CMOS_DrvX_0_SDramEn_5);
    
    \PrState_RNO_0[5]\ : OR2A
      port map(A => \PrState[5]_net_1\, B => SPI_Ok, Y => N_112);
    
    Y_X_WaveEn_RNIGND1 : INV
      port map(A => Y_X_WaveEn_net_1, Y => Y_X_WaveEn_i);
    
    \ACCcnt_RNO_0[5]\ : NOR2B
      port map(A => N_20, B => \ACCcnt[4]_net_1\, Y => N_21);
    
    \PrState_RNO_3[4]\ : OR2B
      port map(A => FrameMk_0_LVDS_ok, B => \PrState[0]_net_1\, Y
         => N_117);
    
    \PrState[7]\ : DFN1P0
      port map(D => CMOS_Ctl_GND, CLK => PLL_Test1_0_Sys_66M_Clk, 
        PRE => PLL_Test1_0_SysRst_O, Q => \PrState[7]_net_1\);
    
    SDramEn_3 : DFN1C0
      port map(D => \PrState_RNI9G29[2]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => CMOS_DrvX_0_SDramEn_3);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \ACCcnt_RNI3P35[2]\ : NOR2
      port map(A => \ACCcnt[2]_net_1\, B => \ACCcnt[3]_net_1\, Y
         => \PrState_ns_0_a3_0_1[7]\);
    
    \ACCcnt_RNO[2]\ : XA1B
      port map(A => \ACCcnt[2]_net_1\, B => N_18, C => 
        \PrState[0]_net_1\, Y => N_128);
    
    \PrState_RNI9G29[2]\ : OR2
      port map(A => \PrState[3]_net_1\, B => \PrState[2]_net_1\, 
        Y => \PrState_RNI9G29[2]_net_1\);
    
    \ACCcnt[4]\ : DFN1E0C0
      port map(D => N_15, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => N_124, Q => \ACCcnt[4]_net_1\);
    
    \PrState[1]\ : DFN1C0
      port map(D => \PrState_RNO[1]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \PrState[1]_net_1\);
    
    \PrState_RNO[5]\ : AO1B
      port map(A => Y_X_WaveOk, B => \PrState[6]_net_1\, C => 
        N_112, Y => \PrState_ns[2]\);
    
    LVDSen_3 : DFN1C0
      port map(D => \PrState[0]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => CMOS_DrvX_0_LVDSen_3);
    
    \PrState_RNO_0[2]\ : OR2B
      port map(A => Y_X_WaveOk, B => \PrState[3]_net_1\, Y => 
        N_120);
    
    \PrState[6]\ : DFN1C0
      port map(D => \PrState_ns[1]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \PrState[6]_net_1\);
    
    LVDSen : DFN1C0
      port map(D => \PrState[0]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => CMOS_DrvX_0_LVDSen);
    
    \PrState_RNO[2]\ : AO1C
      port map(A => Sdram_cmd_0_SDoneFrameOk, B => 
        \PrState[2]_net_1\, C => N_120, Y => \PrState_ns[5]\);
    
    \PrState_RNI5029[1]\ : NOR2
      port map(A => \PrState[1]_net_1\, B => \PrState[0]_net_1\, 
        Y => N_124);
    
    SDramEn_0 : DFN1C0
      port map(D => \PrState_RNI9G29[2]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => CMOS_DrvX_0_SDramEn_0);
    
    SPI_En_0_RNICRT6 : INV
      port map(A => SPI_En_0_net_1, Y => SPI_En_i);
    
    Y_X_WaveEn_RNO : OR2
      port map(A => \PrState[6]_net_1\, B => \PrState[3]_net_1\, 
        Y => \Y_X_WaveEn_RNO\);
    
    \ImageOrQl\ : DFN1P0
      port map(D => \PrState[6]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, PRE => PLL_Test1_0_SysRst_O, Q
         => ImageOrQl);
    
    \ACCcnt[2]\ : DFN1E0C0
      port map(D => N_128, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => N_124, Q => 
        \ACCcnt[2]_net_1\);
    
    \PrState_RNO_0[3]\ : OR2A
      port map(A => \PrState[3]_net_1\, B => Y_X_WaveOk, Y => 
        N_118);
    
    \PrState_RNO[6]\ : AO1A
      port map(A => Y_X_WaveOk, B => \PrState[6]_net_1\, C => 
        \PrState[7]_net_1\, Y => \PrState_ns[1]\);
    
    SDramEn_2 : DFN1C0
      port map(D => \PrState_RNI9G29[2]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => CMOS_DrvX_0_SDramEn_2);
    
    \PrState_RNO[1]\ : NOR2B
      port map(A => Sdram_cmd_0_SDoneFrameOk, B => 
        \PrState[2]_net_1\, Y => \PrState_RNO[1]_net_1\);
    
    \PrState[4]\ : DFN1C0
      port map(D => \PrState_ns[3]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \PrState[4]_net_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \PAT_En\ : DFN1C0
      port map(D => \PrState[4]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => PAT_En);
    
    \ACCcnt_RNIVO35_0[1]\ : NOR2
      port map(A => \ACCcnt[1]_net_1\, B => \ACCcnt[0]_net_1\, Y
         => N_32);
    
    \PrState_RNO_2[4]\ : OR2A
      port map(A => \PrState[4]_net_1\, B => PAT_Ok, Y => N_114);
    
    \PrState[0]\ : DFN1C0
      port map(D => \PrState_ns[7]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \PrState[0]_net_1\);
    
    LVDSen_0 : DFN1C0
      port map(D => \PrState[0]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => CMOS_DrvX_0_LVDSen_0);
    
    SDramEn : DFN1C0
      port map(D => \PrState_RNI9G29[2]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => CMOS_DrvX_0_SDramEn);
    
    \SPI_En_0\ : DFN1C0
      port map(D => \PrState[5]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => SPI_En_0_net_1);
    
    \ACCcnt[3]\ : DFN1E0C0
      port map(D => N_13, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => N_124, Q => \ACCcnt[3]_net_1\);
    
    \SPI_En\ : DFN1C0
      port map(D => \PrState[5]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => SPI_En);
    
    \ACCcnt_RNO[1]\ : NOR3
      port map(A => N_32, B => \PrState[0]_net_1\, C => N_18, Y
         => N_127);
    
    SDramEn_1 : DFN1C0
      port map(D => \PrState_RNI9G29[2]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => CMOS_DrvX_0_SDramEn_1);
    
    \PrState_RNO[3]\ : AO1B
      port map(A => PAT_Ok, B => \PrState[4]_net_1\, C => N_118, 
        Y => \PrState_ns[4]\);
    
    \PrState[3]\ : DFN1C0
      port map(D => \PrState_ns[4]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \PrState[3]_net_1\);
    
    \ACCcnt_RNICDSJ[2]\ : OR3C
      port map(A => N_32, B => \PrState_ns_0_a3_0_1[7]\, C => 
        \PrState_ns_0_a3_0_2[7]\, Y => N_27_i_0);
    
    \ACCcnt_RNO[4]\ : XA1B
      port map(A => \ACCcnt[4]_net_1\, B => N_20, C => 
        \PrState[0]_net_1\, Y => N_15);
    
    \PrState_RNO[0]\ : AO1C
      port map(A => FrameMk_0_LVDS_ok, B => \PrState[0]_net_1\, C
         => N_27_i_0, Y => \PrState_ns[7]\);
    
    \PrState_RNO_0[4]\ : NOR3C
      port map(A => N_115, B => N_114, C => N_117, Y => 
        \PrState_ns_1[3]\);
    
    \ACCcnt_RNO[0]\ : NOR2
      port map(A => \PrState[0]_net_1\, B => \ACCcnt[0]_net_1\, Y
         => ACCcnt_n0);
    
    \Y_X_WaveEn\ : DFN1C0
      port map(D => \Y_X_WaveEn_RNO\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => Y_X_WaveEn_net_1);
    
    \ACCcnt[5]\ : DFN1E0C0
      port map(D => N_17, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => N_124, Q => \ACCcnt[5]_net_1\);
    
    SDramEn_4 : DFN1C0
      port map(D => \PrState_RNI9G29[2]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => CMOS_DrvX_0_SDramEn_4);
    
    \ACCcnt_RNO[3]\ : XA1B
      port map(A => \ACCcnt[3]_net_1\, B => N_19, C => 
        \PrState[0]_net_1\, Y => N_13);
    
    \ACCcnt_RNIGLL7[2]\ : NOR2B
      port map(A => N_18, B => \ACCcnt[2]_net_1\, Y => N_19);
    
    \ACCcnt[0]\ : DFN1E0C0
      port map(D => ACCcnt_n0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => N_124, Q => 
        \ACCcnt[0]_net_1\);
    
    \PrState_RNO_1[4]\ : OR2B
      port map(A => SPI_Ok, B => \PrState[5]_net_1\, Y => N_115);
    
    \PrState_RNO[4]\ : AO1B
      port map(A => \PrState[1]_net_1\, B => N_27_i_0, C => 
        \PrState_ns_1[3]\, Y => \PrState_ns[3]\);
    
    \PrState[5]\ : DFN1C0
      port map(D => \PrState_ns[2]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \PrState[5]_net_1\);
    
    \ACCcnt_RNI2I7A[3]\ : NOR2B
      port map(A => N_19, B => \ACCcnt[3]_net_1\, Y => N_20);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3;
use proasic3.all;

entity SPI_Set is

    port( SPI_En_i                : in    std_logic;
          spi_clock_c             : out   std_logic;
          spi_data_c              : out   std_logic;
          spi_load_c              : out   std_logic;
          SPI_Ok                  : out   std_logic;
          PLL_Test1_0_SysRst_O    : in    std_logic;
          PLL_Test1_0_Sys_66M_Clk : in    std_logic;
          SPI_En                  : in    std_logic;
          SPI_En_0                : in    std_logic
        );

end SPI_Set;

architecture DEF_ARCH of SPI_Set is 

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AOI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component NOR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E0C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AX1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XNOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E0P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

    signal un19_clken_0, \NumCnt[0]_net_1\, \ClkEn\, 
        DivCnt_n1_0_i_0, \DivCnt[0]_net_1\, \DivCnt[1]_net_1\, 
        DivCnt_n1_0_i_a2_1_2, \DivCnt[2]_net_1\, 
        \DivCnt[5]_net_1\, DivCnt_n1_0_i_a2_1_1, 
        \DivCnt[3]_net_1\, \DivCnt[4]_net_1\, N_82, 
        \NumCnt[1]_net_1\, ClkEn_1_sqmuxa_i_0, N_84, N_106, 
        \NumCnt[2]_net_1\, N_86, N_108, \NumCnt[3]_net_1\, N_88, 
        N_137, N_113, N_90, \NumCnt[5]_net_1\, ClkEn_0_sqmuxa_i, 
        N_151, \DivCnt_i[6]\, N_93, N_141, N_103, N_122_i, N_101, 
        N_112, N_99, N_144, N_97, N_107, N_95, N_105, N_312, 
        \PrState[0]_net_1\, \Eof\, N_124, N_126, N_152, N_132, 
        \PrState[1]_net_1\, NumCnt_n0, \NumCnt[4]_net_1\, 
        \ClkEn_RNIGDLA_0\, N_16, \PrState_RNO_2[1]\, \CntEn\, 
        NumCnte, N_156, N_66, \SPI_Shifter[29]_net_1\, N_64, 
        \SPI_Shifter[25]_net_1\, \SPI_Shifter_RNO[23]_net_1\, 
        \SPI_Shifter[24]_net_1\, \SPI_Shifter_RNO[22]_net_1\, 
        \SPI_Shifter[23]_net_1\, \SPI_Shifter_RNO[21]_net_1\, 
        \SPI_Shifter[22]_net_1\, \SPI_Shifter_RNO[20]_net_1\, 
        \SPI_Shifter[21]_net_1\, \SPI_Shifter_RNO[19]_net_1\, 
        \SPI_Shifter[20]_net_1\, \SPI_Shifter_RNO[18]_net_1\, 
        \SPI_Shifter[19]_net_1\, \SPI_Shifter_RNO[17]_net_1\, 
        \SPI_Shifter[18]_net_1\, \SPI_Shifter_RNO[16]_net_1\, 
        \SPI_Shifter[17]_net_1\, \SPI_Shifter_RNO[15]_net_1\, 
        \SPI_Shifter[16]_net_1\, \SPI_Shifter_RNO[14]_net_1\, 
        \SPI_Shifter[15]_net_1\, \SPI_Shifter_RNO[13]_net_1\, 
        \SPI_Shifter[14]_net_1\, \SPI_Shifter_RNO[12]_net_1\, 
        \SPI_Shifter[13]_net_1\, \SPI_Shifter_RNO[11]_net_1\, 
        \SPI_Shifter[12]_net_1\, \SPI_Shifter_RNO[10]_net_1\, 
        \SPI_Shifter[11]_net_1\, \SPI_Shifter_RNO[9]_net_1\, 
        \SPI_Shifter[10]_net_1\, N_32, \SPI_Shifter[9]_net_1\, 
        N_30, \SPI_Shifter[8]_net_1\, N_28, 
        \SPI_Shifter[7]_net_1\, N_26, \SPI_Shifter[6]_net_1\, 
        N_24, \SPI_Shifter[5]_net_1\, N_22, 
        \SPI_Shifter[4]_net_1\, N_20, \SPI_Shifter[3]_net_1\, 
        N_18, \SPI_Shifter[2]_net_1\, N_14, 
        \SPI_Shifter[0]_net_1\, N_12, DivCnt_n0, N_131, 
        \SPI_Shifter[28]_net_1\, N_130, \SPI_Shifter[27]_net_1\, 
        N_129, \SPI_Shifter[26]_net_1\, N_128, 
        \SPI_Shifter[1]_net_1\, \GND\, \VCC\, GND_0, VCC_0
         : std_logic;

begin 


    \SPI_Shifter_RNO[23]\ : NOR2B
      port map(A => SPI_En_0, B => \SPI_Shifter[24]_net_1\, Y => 
        \SPI_Shifter_RNO[23]_net_1\);
    
    \SPI_Shifter[26]\ : DFN1E1C0
      port map(D => N_130, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => \ClkEn_RNIGDLA_0\, Q => 
        \SPI_Shifter[26]_net_1\);
    
    \SPI_Shifter[11]\ : DFN1E1C0
      port map(D => \SPI_Shifter_RNO[11]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => un19_clken_0, Q => \SPI_Shifter[11]_net_1\);
    
    ClkEn_RNIDPR8 : NOR2A
      port map(A => SPI_En_0, B => \ClkEn\, Y => N_124);
    
    \SPI_Shifter[21]\ : DFN1E1C0
      port map(D => \SPI_Shifter_RNO[21]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => un19_clken_0, Q => \SPI_Shifter[21]_net_1\);
    
    \NumCnt_RNO[5]\ : XA1
      port map(A => N_113, B => \NumCnt[5]_net_1\, C => 
        ClkEn_1_sqmuxa_i_0, Y => N_90);
    
    \DivCnt_RNI7QFN1[6]\ : NOR2A
      port map(A => N_151, B => \DivCnt_i[6]\, Y => N_156);
    
    \SPI_Shifter_RNO[19]\ : NOR2B
      port map(A => SPI_En_0, B => \SPI_Shifter[20]_net_1\, Y => 
        \SPI_Shifter_RNO[19]_net_1\);
    
    \NumCnt[2]\ : DFN1E1C0
      port map(D => N_84, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => NumCnte, Q => 
        \NumCnt[2]_net_1\);
    
    \SPI_Shifter_RNO[27]\ : OR2A
      port map(A => SPI_En, B => \SPI_Shifter[28]_net_1\, Y => 
        N_131);
    
    \SPI_Shifter_RNO[11]\ : NOR2B
      port map(A => SPI_En, B => \SPI_Shifter[12]_net_1\, Y => 
        \SPI_Shifter_RNO[11]_net_1\);
    
    \DivCnt_RNO_0[1]\ : NOR3B
      port map(A => DivCnt_n1_0_i_a2_1_1, B => 
        DivCnt_n1_0_i_a2_1_2, C => \DivCnt_i[6]\, Y => N_141);
    
    \DivCnt_RNO[0]\ : NOR2A
      port map(A => ClkEn_1_sqmuxa_i_0, B => \DivCnt[0]_net_1\, Y
         => DivCnt_n0);
    
    \SPI_Shifter_RNO[2]\ : NOR2B
      port map(A => SPI_En, B => \SPI_Shifter[3]_net_1\, Y => 
        N_20);
    
    \SPI_Shifter_RNO[25]\ : OR2A
      port map(A => SPI_En, B => \SPI_Shifter[26]_net_1\, Y => 
        N_129);
    
    \SPI_Shifter_RNO[13]\ : NOR2B
      port map(A => SPI_En, B => \SPI_Shifter[14]_net_1\, Y => 
        \SPI_Shifter_RNO[13]_net_1\);
    
    \SPI_Shifter[13]\ : DFN1E1C0
      port map(D => \SPI_Shifter_RNO[13]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => un19_clken_0, Q => \SPI_Shifter[13]_net_1\);
    
    SPI_Data : DFN1E1C0
      port map(D => N_14, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => un19_clken_0, Q => spi_data_c);
    
    \SPI_Shifter[23]\ : DFN1E1C0
      port map(D => \SPI_Shifter_RNO[23]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => \ClkEn_RNIGDLA_0\, Q => \SPI_Shifter[23]_net_1\);
    
    \NumCnt_RNI7CJ3[1]\ : NOR2B
      port map(A => \NumCnt[1]_net_1\, B => \NumCnt[0]_net_1\, Y
         => N_106);
    
    \NumCnt_RNI1LRA[5]\ : NOR2B
      port map(A => \NumCnt[5]_net_1\, B => N_113, Y => N_152);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \SPI_Ok\ : DFN1C0
      port map(D => \PrState[1]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => SPI_Ok);
    
    \SPI_Shifter_RNO[17]\ : NOR2B
      port map(A => SPI_En_0, B => \SPI_Shifter[18]_net_1\, Y => 
        \SPI_Shifter_RNO[17]_net_1\);
    
    \DivCnt_RNI3OHF1[0]\ : NOR3C
      port map(A => DivCnt_n1_0_i_a2_1_1, B => 
        DivCnt_n1_0_i_a2_1_2, C => \DivCnt[0]_net_1\, Y => N_151);
    
    \SPI_Shifter_RNO[15]\ : NOR2B
      port map(A => SPI_En_0, B => \SPI_Shifter[16]_net_1\, Y => 
        \SPI_Shifter_RNO[15]_net_1\);
    
    \SPI_Shifter[12]\ : DFN1E1C0
      port map(D => \SPI_Shifter_RNO[12]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => un19_clken_0, Q => \SPI_Shifter[12]_net_1\);
    
    \SPI_Shifter_RNO[4]\ : NOR2B
      port map(A => SPI_En, B => \SPI_Shifter[5]_net_1\, Y => 
        N_24);
    
    \SPI_Shifter[22]\ : DFN1E1C0
      port map(D => \SPI_Shifter_RNO[22]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => un19_clken_0, Q => \SPI_Shifter[22]_net_1\);
    
    \SPI_Shifter_RNO[20]\ : NOR2B
      port map(A => SPI_En_0, B => \SPI_Shifter[21]_net_1\, Y => 
        \SPI_Shifter_RNO[20]_net_1\);
    
    ClkEn_RNO : NOR3C
      port map(A => N_151, B => \DivCnt_i[6]\, C => 
        ClkEn_1_sqmuxa_i_0, Y => ClkEn_0_sqmuxa_i);
    
    \SPI_Shifter_RNO[26]\ : OR2A
      port map(A => SPI_En, B => \SPI_Shifter[27]_net_1\, Y => 
        N_130);
    
    \SPI_Shifter[17]\ : DFN1E1C0
      port map(D => \SPI_Shifter_RNO[17]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => un19_clken_0, Q => \SPI_Shifter[17]_net_1\);
    
    \PrState[1]\ : DFN1C0
      port map(D => \PrState_RNO_2[1]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \PrState[1]_net_1\);
    
    \SPI_Shifter_RNO[9]\ : NOR2B
      port map(A => SPI_En, B => \SPI_Shifter[10]_net_1\, Y => 
        \SPI_Shifter_RNO[9]_net_1\);
    
    \SPI_Shifter[27]\ : DFN1E1C0
      port map(D => N_131, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => \ClkEn_RNIGDLA_0\, Q => 
        \SPI_Shifter[27]_net_1\);
    
    \DivCnt_RNIT9ON[2]\ : NOR2B
      port map(A => N_105, B => \DivCnt[2]_net_1\, Y => N_107);
    
    \DivCnt_RNO[3]\ : XA1
      port map(A => \DivCnt[3]_net_1\, B => N_107, C => 
        ClkEn_1_sqmuxa_i_0, Y => N_97);
    
    CntEn : DFN1C0
      port map(D => \PrState[0]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \CntEn\);
    
    SPI_Clock_RNO : NOR2B
      port map(A => SPI_En_0, B => \NumCnt[0]_net_1\, Y => N_16);
    
    \DivCnt[1]\ : DFN1C0
      port map(D => N_93, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \DivCnt[1]_net_1\);
    
    \SPI_Shifter[10]\ : DFN1E1C0
      port map(D => \SPI_Shifter_RNO[10]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => un19_clken_0, Q => \SPI_Shifter[10]_net_1\);
    
    \DivCnt_RNO[6]\ : OR3A
      port map(A => ClkEn_1_sqmuxa_i_0, B => N_151, C => N_122_i, 
        Y => N_103);
    
    \SPI_Shifter_RNO[0]\ : OR2A
      port map(A => SPI_En, B => \SPI_Shifter[1]_net_1\, Y => 
        N_128);
    
    \SPI_Shifter[20]\ : DFN1E1C0
      port map(D => \SPI_Shifter_RNO[20]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => un19_clken_0, Q => \SPI_Shifter[20]_net_1\);
    
    \NumCnt_RNIC8D5[2]\ : NOR2B
      port map(A => \NumCnt[2]_net_1\, B => N_106, Y => N_108);
    
    \DivCnt[6]\ : DFN1P0
      port map(D => N_103, CLK => PLL_Test1_0_Sys_66M_Clk, PRE
         => PLL_Test1_0_SysRst_O, Q => \DivCnt_i[6]\);
    
    \SPI_Shifter_RNO[6]\ : NOR2B
      port map(A => SPI_En, B => \SPI_Shifter[7]_net_1\, Y => 
        N_28);
    
    \SPI_Shifter_RNO[10]\ : NOR2B
      port map(A => SPI_En, B => \SPI_Shifter[11]_net_1\, Y => 
        \SPI_Shifter_RNO[10]_net_1\);
    
    \SPI_Shifter[14]\ : DFN1E1C0
      port map(D => \SPI_Shifter_RNO[14]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => un19_clken_0, Q => \SPI_Shifter[14]_net_1\);
    
    \SPI_Shifter[24]\ : DFN1E1C0
      port map(D => N_64, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => \ClkEn_RNIGDLA_0\, Q => 
        \SPI_Shifter[24]_net_1\);
    
    \NumCnt[1]\ : DFN1E1C0
      port map(D => N_82, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => NumCnte, Q => 
        \NumCnt[1]_net_1\);
    
    \SPI_Shifter_RNO[3]\ : NOR2B
      port map(A => SPI_En, B => \SPI_Shifter[4]_net_1\, Y => 
        N_22);
    
    \SPI_Shifter_RNO[16]\ : NOR2B
      port map(A => SPI_En_0, B => \SPI_Shifter[17]_net_1\, Y => 
        \SPI_Shifter_RNO[16]_net_1\);
    
    \NumCnt_RNO_0[4]\ : AOI1
      port map(A => \NumCnt[3]_net_1\, B => N_108, C => 
        \NumCnt[4]_net_1\, Y => N_137);
    
    \NumCnt_RNO[1]\ : XA1
      port map(A => \NumCnt[0]_net_1\, B => \NumCnt[1]_net_1\, C
         => ClkEn_1_sqmuxa_i_0, Y => N_82);
    
    \DivCnt_RNI2UON[1]\ : NOR3
      port map(A => \DivCnt[2]_net_1\, B => \DivCnt[1]_net_1\, C
         => \DivCnt[5]_net_1\, Y => DivCnt_n1_0_i_a2_1_2);
    
    \DivCnt[3]\ : DFN1C0
      port map(D => N_97, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \DivCnt[3]_net_1\);
    
    \DivCnt[0]\ : DFN1C0
      port map(D => DivCnt_n0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \DivCnt[0]_net_1\);
    
    \NumCnt[5]\ : DFN1E1C0
      port map(D => N_90, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => NumCnte, Q => 
        \NumCnt[5]_net_1\);
    
    \NumCnt[3]\ : DFN1E1C0
      port map(D => N_86, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => NumCnte, Q => 
        \NumCnt[3]_net_1\);
    
    ClkEn_RNIGDLA : AO1C
      port map(A => \NumCnt[0]_net_1\, B => \ClkEn\, C => 
        SPI_En_0, Y => un19_clken_0);
    
    \PrState_RNO[1]\ : OA1
      port map(A => N_312, B => \PrState[1]_net_1\, C => SPI_En_0, 
        Y => \PrState_RNO_2[1]\);
    
    \NumCnt_RNIPC19[4]\ : NOR3C
      port map(A => N_108, B => \NumCnt[3]_net_1\, C => 
        \NumCnt[4]_net_1\, Y => N_113);
    
    Eof_RNIV8J7 : NOR2B
      port map(A => \PrState[0]_net_1\, B => \Eof\, Y => N_312);
    
    \SPI_Shifter_RNO[24]\ : NOR2B
      port map(A => SPI_En_0, B => \SPI_Shifter[25]_net_1\, Y => 
        N_64);
    
    \NumCnt_RNO[0]\ : NOR2A
      port map(A => ClkEn_1_sqmuxa_i_0, B => \NumCnt[0]_net_1\, Y
         => NumCnt_n0);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \DivCnt_RNO[4]\ : NOR3A
      port map(A => ClkEn_1_sqmuxa_i_0, B => N_144, C => N_112, Y
         => N_99);
    
    \DivCnt_RNI3GRF[4]\ : NOR2
      port map(A => \DivCnt[3]_net_1\, B => \DivCnt[4]_net_1\, Y
         => DivCnt_n1_0_i_a2_1_1);
    
    Eof : DFN1E1C0
      port map(D => ClkEn_1_sqmuxa_i_0, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => N_12, Q => \Eof\);
    
    SPI_Clock : DFN1E0C0
      port map(D => N_16, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => N_124, Q => spi_clock_c);
    
    \NumCnt_RNO[3]\ : XA1
      port map(A => N_108, B => \NumCnt[3]_net_1\, C => 
        ClkEn_1_sqmuxa_i_0, Y => N_86);
    
    \NumCnt_RNO[2]\ : XA1
      port map(A => N_106, B => \NumCnt[2]_net_1\, C => 
        ClkEn_1_sqmuxa_i_0, Y => N_84);
    
    \DivCnt_RNO_0[6]\ : AX1C
      port map(A => \DivCnt[5]_net_1\, B => N_112, C => 
        \DivCnt_i[6]\, Y => N_122_i);
    
    \SPI_Shifter_RNO[7]\ : NOR2B
      port map(A => SPI_En, B => \SPI_Shifter[8]_net_1\, Y => 
        N_30);
    
    \DivCnt_RNO[1]\ : NOR3A
      port map(A => ClkEn_1_sqmuxa_i_0, B => N_141, C => 
        DivCnt_n1_0_i_0, Y => N_93);
    
    Eof_RNO : AO1B
      port map(A => N_156, B => N_152, C => ClkEn_1_sqmuxa_i_0, Y
         => N_12);
    
    \DivCnt_RNO[5]\ : XA1
      port map(A => \DivCnt[5]_net_1\, B => N_112, C => 
        ClkEn_1_sqmuxa_i_0, Y => N_101);
    
    \DivCnt_RNI3KC02[6]\ : OR2A
      port map(A => ClkEn_1_sqmuxa_i_0, B => N_156, Y => NumCnte);
    
    ClkEn_RNIGDLA_0 : AO1C
      port map(A => \NumCnt[0]_net_1\, B => \ClkEn\, C => 
        SPI_En_0, Y => \ClkEn_RNIGDLA_0\);
    
    \SPI_Shifter_RNO[5]\ : NOR2B
      port map(A => SPI_En, B => \SPI_Shifter[6]_net_1\, Y => 
        N_26);
    
    \SPI_Shifter[7]\ : DFN1E1C0
      port map(D => N_30, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => \ClkEn_RNIGDLA_0\, Q => 
        \SPI_Shifter[7]_net_1\);
    
    \DivCnt[2]\ : DFN1C0
      port map(D => N_95, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \DivCnt[2]_net_1\);
    
    \PrState[0]\ : DFN1C0
      port map(D => N_132, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \PrState[0]_net_1\);
    
    \SPI_Shifter[0]\ : DFN1E1C0
      port map(D => N_128, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => un19_clken_0, Q => 
        \SPI_Shifter[0]_net_1\);
    
    \SPI_Shifter_RNO[14]\ : NOR2B
      port map(A => SPI_En, B => \SPI_Shifter[15]_net_1\, Y => 
        \SPI_Shifter_RNO[14]_net_1\);
    
    \SPI_Shifter[15]\ : DFN1E1C0
      port map(D => \SPI_Shifter_RNO[15]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => un19_clken_0, Q => \SPI_Shifter[15]_net_1\);
    
    \NumCnt[4]\ : DFN1E1C0
      port map(D => N_88, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => NumCnte, Q => 
        \NumCnt[4]_net_1\);
    
    \SPI_Shifter[25]\ : DFN1E1C0
      port map(D => N_129, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => \ClkEn_RNIGDLA_0\, Q => 
        \SPI_Shifter[25]_net_1\);
    
    \DivCnt_RNITNQF[1]\ : NOR2B
      port map(A => \DivCnt[1]_net_1\, B => \DivCnt[0]_net_1\, Y
         => N_105);
    
    ClkEn : DFN1C0
      port map(D => ClkEn_0_sqmuxa_i, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \ClkEn\);
    
    \SPI_Shifter_RNO[28]\ : NOR2B
      port map(A => SPI_En_0, B => \SPI_Shifter[29]_net_1\, Y => 
        N_66);
    
    \SPI_Shifter[2]\ : DFN1E1C0
      port map(D => N_20, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => \ClkEn_RNIGDLA_0\, Q => 
        \SPI_Shifter[2]_net_1\);
    
    \SPI_Shifter[1]\ : DFN1E1C0
      port map(D => N_18, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => un19_clken_0, Q => 
        \SPI_Shifter[1]_net_1\);
    
    \SPI_Shifter[8]\ : DFN1E1C0
      port map(D => N_32, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => \ClkEn_RNIGDLA_0\, Q => 
        \SPI_Shifter[8]_net_1\);
    
    \NumCnt_RNO[4]\ : NOR3A
      port map(A => ClkEn_1_sqmuxa_i_0, B => N_137, C => N_113, Y
         => N_88);
    
    \DivCnt_RNI0QJ71[4]\ : NOR3C
      port map(A => \DivCnt[3]_net_1\, B => N_107, C => 
        \DivCnt[4]_net_1\, Y => N_112);
    
    \DivCnt[5]\ : DFN1C0
      port map(D => N_101, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \DivCnt[5]_net_1\);
    
    \SPI_Shifter_RNO[22]\ : NOR2B
      port map(A => SPI_En_0, B => \SPI_Shifter[23]_net_1\, Y => 
        \SPI_Shifter_RNO[22]_net_1\);
    
    \SPI_Shifter[6]\ : DFN1E1C0
      port map(D => N_28, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => \ClkEn_RNIGDLA_0\, Q => 
        \SPI_Shifter[6]_net_1\);
    
    \SPI_Shifter[4]\ : DFN1E1C0
      port map(D => N_24, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => \ClkEn_RNIGDLA_0\, Q => 
        \SPI_Shifter[4]_net_1\);
    
    \SPI_Shifter[19]\ : DFN1E1C0
      port map(D => \SPI_Shifter_RNO[19]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => un19_clken_0, Q => \SPI_Shifter[19]_net_1\);
    
    SPI_Load_RNO : OR2B
      port map(A => SPI_En_0, B => N_152, Y => N_126);
    
    \SPI_Shifter[29]\ : DFN1E1C0
      port map(D => SPI_En_i, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => \ClkEn_RNIGDLA_0\, Q => 
        \SPI_Shifter[29]_net_1\);
    
    \SPI_Shifter[9]\ : DFN1E1C0
      port map(D => \SPI_Shifter_RNO[9]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => \ClkEn_RNIGDLA_0\, Q => \SPI_Shifter[9]_net_1\);
    
    \DivCnt_RNO_1[1]\ : XNOR2
      port map(A => \DivCnt[0]_net_1\, B => \DivCnt[1]_net_1\, Y
         => DivCnt_n1_0_i_0);
    
    \SPI_Shifter_RNO[1]\ : NOR2B
      port map(A => SPI_En, B => \SPI_Shifter[2]_net_1\, Y => 
        N_18);
    
    \PrState_RNO[0]\ : NOR3A
      port map(A => SPI_En_0, B => N_312, C => \PrState[1]_net_1\, 
        Y => N_132);
    
    \DivCnt_RNO_0[4]\ : AOI1
      port map(A => N_107, B => \DivCnt[3]_net_1\, C => 
        \DivCnt[4]_net_1\, Y => N_144);
    
    \SPI_Shifter_RNO[8]\ : NOR2B
      port map(A => SPI_En, B => \SPI_Shifter[9]_net_1\, Y => 
        N_32);
    
    \SPI_Shifter_RNO[18]\ : NOR2B
      port map(A => SPI_En_0, B => \SPI_Shifter[19]_net_1\, Y => 
        \SPI_Shifter_RNO[18]_net_1\);
    
    CntEn_RNISPS8 : NOR2B
      port map(A => SPI_En_0, B => \CntEn\, Y => 
        ClkEn_1_sqmuxa_i_0);
    
    SPI_Data_RNO : NOR2B
      port map(A => SPI_En, B => \SPI_Shifter[0]_net_1\, Y => 
        N_14);
    
    \SPI_Shifter[18]\ : DFN1E1C0
      port map(D => \SPI_Shifter_RNO[18]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => un19_clken_0, Q => \SPI_Shifter[18]_net_1\);
    
    \SPI_Shifter[5]\ : DFN1E1C0
      port map(D => N_26, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => \ClkEn_RNIGDLA_0\, Q => 
        \SPI_Shifter[5]_net_1\);
    
    \SPI_Shifter[28]\ : DFN1E1C0
      port map(D => N_66, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => \ClkEn_RNIGDLA_0\, Q => 
        \SPI_Shifter[28]_net_1\);
    
    \DivCnt_RNO[2]\ : XA1
      port map(A => \DivCnt[2]_net_1\, B => N_105, C => 
        ClkEn_1_sqmuxa_i_0, Y => N_95);
    
    \DivCnt[4]\ : DFN1C0
      port map(D => N_99, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \DivCnt[4]_net_1\);
    
    \SPI_Shifter_RNO[12]\ : NOR2B
      port map(A => SPI_En, B => \SPI_Shifter[13]_net_1\, Y => 
        \SPI_Shifter_RNO[12]_net_1\);
    
    \SPI_Shifter_RNO[21]\ : NOR2B
      port map(A => SPI_En_0, B => \SPI_Shifter[22]_net_1\, Y => 
        \SPI_Shifter_RNO[21]_net_1\);
    
    \SPI_Shifter[3]\ : DFN1E1C0
      port map(D => N_22, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => \ClkEn_RNIGDLA_0\, Q => 
        \SPI_Shifter[3]_net_1\);
    
    SPI_Load : DFN1E0P0
      port map(D => N_126, CLK => PLL_Test1_0_Sys_66M_Clk, PRE
         => PLL_Test1_0_SysRst_O, E => N_124, Q => spi_load_c);
    
    \NumCnt[0]\ : DFN1E1C0
      port map(D => NumCnt_n0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => NumCnte, Q => 
        \NumCnt[0]_net_1\);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    \SPI_Shifter[16]\ : DFN1E1C0
      port map(D => \SPI_Shifter_RNO[16]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => un19_clken_0, Q => \SPI_Shifter[16]_net_1\);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3;
use proasic3.all;

entity PixelArrayTiming is

    port( PAT_Ok                  : out   std_logic;
          mem_HL_c                : out   std_logic;
          precharge_c             : out   std_logic;
          CMOS_sample_c           : out   std_logic;
          CMOS_reset_c            : out   std_logic;
          PAT_En                  : in    std_logic;
          PLL_Test1_0_SysRst_O    : in    std_logic;
          PLL_Test1_0_Sys_66M_Clk : in    std_logic
        );

end PixelArrayTiming;

architecture DEF_ARCH of PixelArrayTiming is 

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OAI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component AO1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E0P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component NOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1D
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XAI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \ClkEn_1\, ClkEn_4, \ClkEn_0\, DivCnt_n6_0_i_0, N_41, 
        \DivCnt[0]_net_1\, \InitCnt_5_i_a3_1[0]\, 
        \InitCnt[0]_net_1\, un1_initcnt14_i_a3_0, 
        un27_clken_0_o2_0, un27_clken_0_a2_0, N_47, N_80, 
        un1_pat_en_1_0_a2_0, \InitCnt[1]_net_1\, 
        \InitCnt[4]_net_1\, un27_clken_0_a2_0_9, 
        un27_clken_0_a2_0_6, \InitCnt[15]_net_1\, 
        \InitCnt[14]_net_1\, un27_clken_0_a2_0_8, 
        un27_clken_0_a2_0_4, \InitCnt[11]_net_1\, 
        \InitCnt[10]_net_1\, un27_clken_0_a2_0_7, 
        un27_clken_0_a2_0_2, \InitCnt[7]_net_1\, 
        \InitCnt[6]_net_1\, \InitCnt[5]_net_1\, 
        \InitCnt[17]_net_1\, \InitCnt[16]_net_1\, 
        \InitCnt[12]_net_1\, \InitCnt[13]_net_1\, 
        \InitCnt[8]_net_1\, \InitCnt[9]_net_1\, ClkEn_4_0_a4_0, 
        \DivCnt[6]_net_1\, DivCnt_n1_0_i_1, \DivCnt[1]_net_1\, 
        DivCnt_n1_0_i_a2_2, \DivCnt[2]_net_1\, \DivCnt[5]_net_1\, 
        \DivCnt[4]_net_1\, \DivCnt[3]_net_1\, N_8, N_17, N_10, 
        N_18, N_12, N_19, N_14, N_20, N_94, N_6, N_16, N_171, 
        N_69, N_82, \InitCnt[3]_net_1\, N_49, N_73, N_180, 
        \InitCnt_RNO[5]_net_1\, I_63, \InitCnt_RNO[3]_net_1\, 
        I_72, N_44, I_67, N_46, I_73, \InitCnt_RNO[8]_net_1\, 
        I_69, \InitCnt_RNO[6]_net_1\, I_65, 
        \InitCnt_RNO[4]_net_1\, I_61, \InitCnt_RNO[2]_net_1\, 
        I_68, \InitCnt_RNO[1]_net_1\, I_62, 
        \InitCnt_RNO[17]_net_1\, I_74, \InitCnt_RNO[14]_net_1\, 
        I_64, \InitCnt_RNO[13]_net_1\, I_58, 
        \InitCnt_RNO[9]_net_1\, I_70, \InitCnt_RNO[16]_net_1\, 
        I_71, \InitCnt_RNO[15]_net_1\, I_66, 
        \InitCnt_RNO[12]_net_1\, I_59, \InitCnt_RNO[11]_net_1\, 
        I_57, \InitCnt[2]_net_1\, N_48, N_78, N_40, 
        \DWACT_ADD_CI_0_partial_sum[0]\, un1_pat_en_1, un52_clken, 
        un39_clken, un27_clken, N_68, DivCnt_n0, \ClkEn\, 
        \DWACT_ADD_CI_0_pog_array_1_6[0]\, 
        \DWACT_ADD_CI_0_pog_array_0_13[0]\, 
        \DWACT_ADD_CI_0_pog_array_0_14[0]\, 
        \DWACT_ADD_CI_0_pog_array_2_1[0]\, 
        \DWACT_ADD_CI_0_pog_array_1_3[0]\, 
        \DWACT_ADD_CI_0_pog_array_1_4[0]\, 
        \DWACT_ADD_CI_0_pog_array_2_2[0]\, 
        \DWACT_ADD_CI_0_pog_array_1_5[0]\, 
        \DWACT_ADD_CI_0_pog_array_0_11[0]\, 
        \DWACT_ADD_CI_0_pog_array_0_12[0]\, 
        \DWACT_ADD_CI_0_pog_array_1_2[0]\, 
        \DWACT_ADD_CI_0_pog_array_0_5[0]\, 
        \DWACT_ADD_CI_0_pog_array_0_6[0]\, 
        \DWACT_ADD_CI_0_pog_array_0_9[0]\, 
        \DWACT_ADD_CI_0_pog_array_0_10[0]\, 
        \DWACT_ADD_CI_0_pog_array_1_1[0]\, 
        \DWACT_ADD_CI_0_pog_array_0_3[0]\, 
        \DWACT_ADD_CI_0_pog_array_0_4[0]\, 
        \DWACT_ADD_CI_0_pog_array_2[0]\, 
        \DWACT_ADD_CI_0_pog_array_0_7[0]\, 
        \DWACT_ADD_CI_0_pog_array_0_8[0]\, 
        \DWACT_ADD_CI_0_pog_array_1[0]\, 
        \DWACT_ADD_CI_0_pog_array_0_1[0]\, 
        \DWACT_ADD_CI_0_pog_array_0_2[0]\, 
        \DWACT_ADD_CI_0_pog_array_3[0]\, 
        \DWACT_ADD_CI_0_g_array_12_7[0]\, 
        \DWACT_ADD_CI_0_pog_array_0_15[0]\, 
        \DWACT_ADD_CI_0_g_array_4[0]\, 
        \DWACT_ADD_CI_0_g_array_0_16[0]\, 
        \DWACT_ADD_CI_0_g_array_11_2[0]\, 
        \DWACT_ADD_CI_0_g_array_10[0]\, 
        \DWACT_ADD_CI_0_g_array_1_6[0]\, 
        \DWACT_ADD_CI_0_g_array_12[0]\, 
        \DWACT_ADD_CI_0_g_array_1[0]\, 
        \DWACT_ADD_CI_0_g_array_0_2[0]\, 
        \DWACT_ADD_CI_0_g_array_12_5[0]\, 
        \DWACT_ADD_CI_0_g_array_0_12[0]\, 
        \DWACT_ADD_CI_0_g_array_11[0]\, 
        \DWACT_ADD_CI_0_g_array_2[0]\, 
        \DWACT_ADD_CI_0_g_array_1_2[0]\, 
        \DWACT_ADD_CI_0_g_array_2_1[0]\, 
        \DWACT_ADD_CI_0_g_array_1_3[0]\, 
        \DWACT_ADD_CI_0_g_array_12_4[0]\, 
        \DWACT_ADD_CI_0_g_array_11_1[0]\, 
        \DWACT_ADD_CI_0_g_array_0_10[0]\, 
        \DWACT_ADD_CI_0_g_array_1_1[0]\, 
        \DWACT_ADD_CI_0_g_array_3[0]\, 
        \DWACT_ADD_CI_0_g_array_3_1[0]\, 
        \DWACT_ADD_CI_0_g_array_12_3[0]\, 
        \DWACT_ADD_CI_0_g_array_0_8[0]\, 
        \DWACT_ADD_CI_0_g_array_12_2[0]\, 
        \DWACT_ADD_CI_0_g_array_0_6[0]\, 
        \DWACT_ADD_CI_0_g_array_2_2[0]\, 
        \DWACT_ADD_CI_0_g_array_2_3[0]\, 
        \DWACT_ADD_CI_0_g_array_12_1[0]\, 
        \DWACT_ADD_CI_0_g_array_0_4[0]\, 
        \DWACT_ADD_CI_0_g_array_1_4[0]\, 
        \DWACT_ADD_CI_0_g_array_1_5[0]\, 
        \DWACT_ADD_CI_0_g_array_1_7[0]\, 
        \DWACT_ADD_CI_0_g_array_0_14[0]\, 
        \DWACT_ADD_CI_0_g_array_0_15[0]\, 
        \DWACT_ADD_CI_0_g_array_12_6[0]\, 
        \DWACT_ADD_CI_0_g_array_0_7[0]\, 
        \DWACT_ADD_CI_0_g_array_0_13[0]\, 
        \DWACT_ADD_CI_0_g_array_0_5[0]\, 
        \DWACT_ADD_CI_0_g_array_0_11[0]\, 
        \DWACT_ADD_CI_0_g_array_0_3[0]\, 
        \DWACT_ADD_CI_0_g_array_0_9[0]\, 
        \DWACT_ADD_CI_0_pog_array_0[0]\, \DWACT_ADD_CI_0_TMP[0]\, 
        \DWACT_ADD_CI_0_g_array_0_1[0]\, 
        \DWACT_ADD_CI_0_partial_sum[17]\, 
        \DWACT_ADD_CI_0_partial_sum[10]\, 
        \DWACT_ADD_CI_0_partial_sum[3]\, 
        \DWACT_ADD_CI_0_partial_sum[16]\, 
        \DWACT_ADD_CI_0_partial_sum[9]\, 
        \DWACT_ADD_CI_0_partial_sum[8]\, 
        \DWACT_ADD_CI_0_partial_sum[2]\, 
        \DWACT_ADD_CI_0_partial_sum[7]\, 
        \DWACT_ADD_CI_0_partial_sum[15]\, 
        \DWACT_ADD_CI_0_partial_sum[6]\, 
        \DWACT_ADD_CI_0_partial_sum[14]\, 
        \DWACT_ADD_CI_0_partial_sum[5]\, 
        \DWACT_ADD_CI_0_partial_sum[1]\, 
        \DWACT_ADD_CI_0_partial_sum[4]\, 
        \DWACT_ADD_CI_0_partial_sum[12]\, 
        \DWACT_ADD_CI_0_partial_sum[13]\, 
        \DWACT_ADD_CI_0_partial_sum[11]\, \GND\, \VCC\, GND_0, 
        VCC_0 : std_logic;

begin 


    \DivCnt_RNITNF91[0]\ : NOR3C
      port map(A => \DivCnt[0]_net_1\, B => N_41, C => 
        ClkEn_4_0_a4_0, Y => ClkEn_4);
    
    un1_InitCnt_I_108 : AND2
      port map(A => \DWACT_ADD_CI_0_pog_array_0_3[0]\, B => 
        \DWACT_ADD_CI_0_pog_array_0_4[0]\, Y => 
        \DWACT_ADD_CI_0_pog_array_1_1[0]\);
    
    ClkEn_1 : DFN1C0
      port map(D => ClkEn_4, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \ClkEn_1\);
    
    un1_InitCnt_I_83 : AO1
      port map(A => \DWACT_ADD_CI_0_pog_array_2[0]\, B => 
        \DWACT_ADD_CI_0_g_array_2[0]\, C => 
        \DWACT_ADD_CI_0_g_array_2_1[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_3[0]\);
    
    un1_InitCnt_I_51 : XOR2
      port map(A => \InitCnt[15]_net_1\, B => \ClkEn\, Y => 
        \DWACT_ADD_CI_0_partial_sum[15]\);
    
    \InitCnt[2]\ : DFN1C0
      port map(D => \InitCnt_RNO[2]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \InitCnt[2]_net_1\);
    
    \InitCnt[0]\ : DFN1C0
      port map(D => N_40, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \InitCnt[0]_net_1\);
    
    un1_InitCnt_I_33 : XOR2
      port map(A => \InitCnt[11]_net_1\, B => \ClkEn_1\, Y => 
        \DWACT_ADD_CI_0_pog_array_0_10[0]\);
    
    \InitCnt[5]\ : DFN1C0
      port map(D => \InitCnt_RNO[5]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \InitCnt[5]_net_1\);
    
    un1_InitCnt_I_69 : XOR2
      port map(A => \DWACT_ADD_CI_0_partial_sum[8]\, B => 
        \DWACT_ADD_CI_0_g_array_3[0]\, Y => I_69);
    
    un1_InitCnt_I_67 : XOR2
      port map(A => \DWACT_ADD_CI_0_partial_sum[7]\, B => 
        \DWACT_ADD_CI_0_g_array_12_2[0]\, Y => I_67);
    
    un1_InitCnt_I_73 : XOR2
      port map(A => \DWACT_ADD_CI_0_partial_sum[10]\, B => 
        \DWACT_ADD_CI_0_g_array_11_1[0]\, Y => I_73);
    
    \InitCnt_RNI1U26[0]\ : OR2A
      port map(A => \ClkEn_0\, B => \InitCnt[0]_net_1\, Y => 
        un1_initcnt14_i_a3_0);
    
    \InitCnt_RNO[10]\ : OA1A
      port map(A => PAT_En, B => I_73, C => N_73, Y => N_46);
    
    un1_InitCnt_I_64 : XOR2
      port map(A => \DWACT_ADD_CI_0_partial_sum[14]\, B => 
        \DWACT_ADD_CI_0_g_array_11_2[0]\, Y => I_64);
    
    \PAT_Ok\ : DFN1E1C0
      port map(D => PAT_En, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => N_180, Q => PAT_Ok);
    
    \InitCnt_RNO[16]\ : NOR2A
      port map(A => I_71, B => N_180, Y => 
        \InitCnt_RNO[16]_net_1\);
    
    sample_RNO : OR2B
      port map(A => N_94, B => N_48, Y => un52_clken);
    
    \InitCnt_RNIVNPD2[0]\ : OR3B
      port map(A => N_94, B => un1_pat_en_1_0_a2_0, C => 
        \InitCnt_5_i_a3_1[0]\, Y => N_73);
    
    \InitCnt[13]\ : DFN1C0
      port map(D => \InitCnt_RNO[13]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \InitCnt[13]_net_1\);
    
    \DivCnt[0]\ : DFN1C0
      port map(D => DivCnt_n0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \DivCnt[0]_net_1\);
    
    precharge_RNO_1 : OR2
      port map(A => \InitCnt[2]_net_1\, B => \InitCnt[1]_net_1\, 
        Y => N_49);
    
    un1_InitCnt_I_114 : AND2
      port map(A => \DWACT_ADD_CI_0_pog_array_0_13[0]\, B => 
        \DWACT_ADD_CI_0_pog_array_0_14[0]\, Y => 
        \DWACT_ADD_CI_0_pog_array_1_6[0]\);
    
    \DivCnt_RNITOAF[2]\ : NOR2B
      port map(A => N_17, B => \DivCnt[2]_net_1\, Y => N_18);
    
    un1_InitCnt_I_112 : AND2
      port map(A => \DWACT_ADD_CI_0_pog_array_1_5[0]\, B => 
        \DWACT_ADD_CI_0_pog_array_1_6[0]\, Y => 
        \DWACT_ADD_CI_0_pog_array_2_2[0]\);
    
    \InitCnt_RNIVNPD2_0[0]\ : OR2B
      port map(A => PAT_En, B => N_69, Y => N_180);
    
    \InitCnt_RNI4RMD[4]\ : AO1A
      port map(A => \InitCnt[4]_net_1\, B => N_47, C => N_78, Y
         => N_48);
    
    un1_InitCnt_I_13 : AND2
      port map(A => \InitCnt[9]_net_1\, B => \ClkEn_0\, Y => 
        \DWACT_ADD_CI_0_g_array_0_9[0]\);
    
    un1_InitCnt_I_65 : XOR2
      port map(A => \DWACT_ADD_CI_0_partial_sum[6]\, B => 
        \DWACT_ADD_CI_0_g_array_11[0]\, Y => I_65);
    
    un1_InitCnt_I_110 : AND2
      port map(A => \DWACT_ADD_CI_0_pog_array_0_5[0]\, B => 
        \DWACT_ADD_CI_0_pog_array_0_6[0]\, Y => 
        \DWACT_ADD_CI_0_pog_array_1_2[0]\);
    
    un1_InitCnt_I_66 : XOR2
      port map(A => \DWACT_ADD_CI_0_partial_sum[15]\, B => 
        \DWACT_ADD_CI_0_g_array_12_6[0]\, Y => I_66);
    
    un1_InitCnt_I_62 : XOR2
      port map(A => \DWACT_ADD_CI_0_partial_sum[1]\, B => 
        \DWACT_ADD_CI_0_TMP[0]\, Y => I_62);
    
    \DivCnt[5]\ : DFN1C0
      port map(D => N_14, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \DivCnt[5]_net_1\);
    
    un1_InitCnt_I_9 : AND2
      port map(A => \InitCnt[3]_net_1\, B => \ClkEn\, Y => 
        \DWACT_ADD_CI_0_g_array_0_3[0]\);
    
    \DivCnt_RNO[2]\ : XA1
      port map(A => \DivCnt[2]_net_1\, B => N_17, C => PAT_En, Y
         => N_8);
    
    \DivCnt_RNO[1]\ : AOI1
      port map(A => N_41, B => \DivCnt[6]_net_1\, C => 
        DivCnt_n1_0_i_1, Y => N_6);
    
    \InitCnt[4]\ : DFN1C0
      port map(D => \InitCnt_RNO[4]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \InitCnt[4]_net_1\);
    
    mem_HL_RNO : OAI1
      port map(A => N_48, B => un27_clken_0_o2_0, C => N_94, Y
         => un27_clken);
    
    \InitCnt_RNIVQU3[8]\ : NOR2
      port map(A => \InitCnt[8]_net_1\, B => \InitCnt[9]_net_1\, 
        Y => un27_clken_0_a2_0_2);
    
    ClkEn : DFN1C0
      port map(D => ClkEn_4, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \ClkEn\);
    
    \InitCnt_RNO[0]\ : OA1A
      port map(A => PAT_En, B => \DWACT_ADD_CI_0_partial_sum[0]\, 
        C => N_73, Y => N_40);
    
    \InitCnt[8]\ : DFN1C0
      port map(D => \InitCnt_RNO[8]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \InitCnt[8]_net_1\);
    
    \InitCnt_RNI2I5Q1[6]\ : NOR3C
      port map(A => un27_clken_0_a2_0_8, B => un27_clken_0_a2_0_7, 
        C => un27_clken_0_a2_0_9, Y => N_94);
    
    sample : DFN1E1P0
      port map(D => un52_clken, CLK => PLL_Test1_0_Sys_66M_Clk, 
        PRE => PLL_Test1_0_SysRst_O, E => \ClkEn_0\, Q => 
        CMOS_sample_c);
    
    un1_InitCnt_I_50 : XOR2
      port map(A => \InitCnt[3]_net_1\, B => \ClkEn\, Y => 
        \DWACT_ADD_CI_0_partial_sum[3]\);
    
    \InitCnt_RNO[4]\ : NOR2A
      port map(A => I_61, B => N_180, Y => \InitCnt_RNO[4]_net_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \DivCnt_RNI0VHP[4]\ : NOR2B
      port map(A => N_19, B => \DivCnt[4]_net_1\, Y => N_20);
    
    \InitCnt_RNO[11]\ : NOR2A
      port map(A => I_57, B => N_180, Y => 
        \InitCnt_RNO[11]_net_1\);
    
    \DivCnt_RNIUBEK[3]\ : NOR2B
      port map(A => N_18, B => \DivCnt[3]_net_1\, Y => N_19);
    
    \InitCnt_RNO[2]\ : NOR2A
      port map(A => I_68, B => N_180, Y => \InitCnt_RNO[2]_net_1\);
    
    un1_InitCnt_I_59 : XOR2
      port map(A => \DWACT_ADD_CI_0_partial_sum[12]\, B => 
        \DWACT_ADD_CI_0_g_array_10[0]\, Y => I_59);
    
    \DivCnt_RNO_1[6]\ : AO1B
      port map(A => N_41, B => \DivCnt[0]_net_1\, C => PAT_En, Y
         => DivCnt_n6_0_i_0);
    
    reset : DFN1E0P0
      port map(D => un1_pat_en_1, CLK => PLL_Test1_0_Sys_66M_Clk, 
        PRE => PLL_Test1_0_SysRst_O, E => N_68, Q => CMOS_reset_c);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    un1_InitCnt_I_57 : XOR2
      port map(A => \DWACT_ADD_CI_0_partial_sum[11]\, B => 
        \DWACT_ADD_CI_0_g_array_12_4[0]\, Y => I_57);
    
    \InitCnt[6]\ : DFN1C0
      port map(D => \InitCnt_RNO[6]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \InitCnt[6]_net_1\);
    
    un1_InitCnt_I_109 : AND2
      port map(A => \DWACT_ADD_CI_0_pog_array_0_9[0]\, B => 
        \DWACT_ADD_CI_0_pog_array_0_10[0]\, Y => 
        \DWACT_ADD_CI_0_pog_array_1_4[0]\);
    
    un1_InitCnt_I_54 : XOR2
      port map(A => \InitCnt[14]_net_1\, B => \ClkEn\, Y => 
        \DWACT_ADD_CI_0_partial_sum[14]\);
    
    un1_InitCnt_I_7 : AND2
      port map(A => \InitCnt[16]_net_1\, B => \ClkEn\, Y => 
        \DWACT_ADD_CI_0_g_array_0_16[0]\);
    
    un1_InitCnt_I_104 : AND2
      port map(A => \DWACT_ADD_CI_0_pog_array_2_1[0]\, B => 
        \DWACT_ADD_CI_0_pog_array_2_2[0]\, Y => 
        \DWACT_ADD_CI_0_pog_array_3[0]\);
    
    \DivCnt_RNI2PAF[1]\ : NOR3
      port map(A => \DivCnt[2]_net_1\, B => \DivCnt[1]_net_1\, C
         => \DivCnt[5]_net_1\, Y => DivCnt_n1_0_i_a2_2);
    
    un1_InitCnt_I_98 : AO1
      port map(A => \DWACT_ADD_CI_0_pog_array_1_2[0]\, B => 
        \DWACT_ADD_CI_0_g_array_1_2[0]\, C => 
        \DWACT_ADD_CI_0_g_array_1_3[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_2_1[0]\);
    
    un1_InitCnt_I_102 : AO1
      port map(A => \DWACT_ADD_CI_0_pog_array_1_5[0]\, B => 
        \DWACT_ADD_CI_0_g_array_10[0]\, C => 
        \DWACT_ADD_CI_0_g_array_1_6[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_11_2[0]\);
    
    un1_InitCnt_I_48 : XOR2
      port map(A => \InitCnt[16]_net_1\, B => \ClkEn\, Y => 
        \DWACT_ADD_CI_0_partial_sum[16]\);
    
    reset_RNO_0 : NOR2A
      port map(A => PAT_En, B => \ClkEn_0\, Y => N_68);
    
    un1_InitCnt_I_63 : XOR2
      port map(A => \DWACT_ADD_CI_0_partial_sum[5]\, B => 
        \DWACT_ADD_CI_0_g_array_12_1[0]\, Y => I_63);
    
    un1_InitCnt_I_91 : AO1
      port map(A => \DWACT_ADD_CI_0_pog_array_2_2[0]\, B => 
        \DWACT_ADD_CI_0_g_array_2_2[0]\, C => 
        \DWACT_ADD_CI_0_g_array_2_3[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_3_1[0]\);
    
    un1_InitCnt_I_41 : XOR2
      port map(A => \InitCnt[4]_net_1\, B => \ClkEn_1\, Y => 
        \DWACT_ADD_CI_0_partial_sum[4]\);
    
    \InitCnt[11]\ : DFN1C0
      port map(D => \InitCnt_RNO[11]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \InitCnt[11]_net_1\);
    
    un1_InitCnt_I_55 : XOR2
      port map(A => \InitCnt[9]_net_1\, B => \ClkEn\, Y => 
        \DWACT_ADD_CI_0_partial_sum[9]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    un1_InitCnt_I_100 : AO1
      port map(A => \DWACT_ADD_CI_0_pog_array_0_11[0]\, B => 
        \DWACT_ADD_CI_0_g_array_10[0]\, C => 
        \DWACT_ADD_CI_0_g_array_0_12[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_12_5[0]\);
    
    un1_InitCnt_I_56 : XOR2
      port map(A => \InitCnt[6]_net_1\, B => \ClkEn\, Y => 
        \DWACT_ADD_CI_0_partial_sum[6]\);
    
    un1_InitCnt_I_28 : XOR2
      port map(A => \InitCnt[14]_net_1\, B => \ClkEn_1\, Y => 
        \DWACT_ADD_CI_0_pog_array_0_13[0]\);
    
    un1_InitCnt_I_52 : XOR2
      port map(A => \InitCnt[10]_net_1\, B => \ClkEn\, Y => 
        \DWACT_ADD_CI_0_partial_sum[10]\);
    
    \DivCnt[1]\ : DFN1C0
      port map(D => N_6, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \DivCnt[1]_net_1\);
    
    un1_InitCnt_I_1 : AND2
      port map(A => \InitCnt[0]_net_1\, B => \ClkEn_0\, Y => 
        \DWACT_ADD_CI_0_TMP[0]\);
    
    un1_InitCnt_I_21 : AND2
      port map(A => \InitCnt[5]_net_1\, B => \ClkEn_0\, Y => 
        \DWACT_ADD_CI_0_g_array_0_5[0]\);
    
    precharge_RNO : OAI1
      port map(A => N_78, B => N_82, C => N_94, Y => un39_clken);
    
    \InitCnt_RNIJAT3[2]\ : OR2
      port map(A => \InitCnt[3]_net_1\, B => \InitCnt[2]_net_1\, 
        Y => N_47);
    
    \InitCnt[17]\ : DFN1C0
      port map(D => \InitCnt_RNO[17]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \InitCnt[17]_net_1\);
    
    un1_InitCnt_I_113 : AND2
      port map(A => \DWACT_ADD_CI_0_pog_array_1_3[0]\, B => 
        \DWACT_ADD_CI_0_pog_array_1_4[0]\, Y => 
        \DWACT_ADD_CI_0_pog_array_2_1[0]\);
    
    un1_InitCnt_I_88 : AO1
      port map(A => \DWACT_ADD_CI_0_pog_array_0_14[0]\, B => 
        \DWACT_ADD_CI_0_g_array_0_14[0]\, C => 
        \DWACT_ADD_CI_0_g_array_0_15[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_1_7[0]\);
    
    \DivCnt[4]\ : DFN1C0
      port map(D => N_12, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \DivCnt[4]_net_1\);
    
    un1_InitCnt_I_81 : AO1
      port map(A => \DWACT_ADD_CI_0_pog_array_0_4[0]\, B => 
        \DWACT_ADD_CI_0_g_array_0_4[0]\, C => 
        \DWACT_ADD_CI_0_g_array_0_5[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_1_2[0]\);
    
    un1_InitCnt_I_78 : AO1
      port map(A => \DWACT_ADD_CI_0_pog_array_2_1[0]\, B => 
        \DWACT_ADD_CI_0_g_array_3[0]\, C => 
        \DWACT_ADD_CI_0_g_array_2_2[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_10[0]\);
    
    un1_InitCnt_I_31 : XOR2
      port map(A => \InitCnt[5]_net_1\, B => \ClkEn_1\, Y => 
        \DWACT_ADD_CI_0_pog_array_0_4[0]\);
    
    \InitCnt_RNI6LQ7[1]\ : NOR3A
      port map(A => \InitCnt[4]_net_1\, B => \InitCnt[1]_net_1\, 
        C => N_47, Y => N_78);
    
    un1_InitCnt_I_71 : XOR2
      port map(A => \DWACT_ADD_CI_0_partial_sum[16]\, B => 
        \DWACT_ADD_CI_0_g_array_4[0]\, Y => I_71);
    
    \InitCnt_RNO[12]\ : NOR2A
      port map(A => I_59, B => N_180, Y => 
        \InitCnt_RNO[12]_net_1\);
    
    \InitCnt[15]\ : DFN1C0
      port map(D => \InitCnt_RNO[15]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \InitCnt[15]_net_1\);
    
    precharge_RNO_0 : NOR3B
      port map(A => \InitCnt[3]_net_1\, B => N_49, C => 
        \InitCnt[4]_net_1\, Y => N_82);
    
    \DivCnt_RNO[4]\ : XA1
      port map(A => \DivCnt[4]_net_1\, B => N_19, C => PAT_En, Y
         => N_12);
    
    un1_InitCnt_I_107 : AND2
      port map(A => \DWACT_ADD_CI_0_pog_array_1_1[0]\, B => 
        \DWACT_ADD_CI_0_pog_array_1_2[0]\, Y => 
        \DWACT_ADD_CI_0_pog_array_2[0]\);
    
    \InitCnt[10]\ : DFN1C0
      port map(D => N_46, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \InitCnt[10]_net_1\);
    
    \InitCnt[1]\ : DFN1C0
      port map(D => \InitCnt_RNO[1]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \InitCnt[1]_net_1\);
    
    un1_InitCnt_I_111 : AND2
      port map(A => \DWACT_ADD_CI_0_pog_array_0_11[0]\, B => 
        \DWACT_ADD_CI_0_pog_array_0_12[0]\, Y => 
        \DWACT_ADD_CI_0_pog_array_1_5[0]\);
    
    un1_InitCnt_I_18 : AND2
      port map(A => \InitCnt[1]_net_1\, B => \ClkEn_0\, Y => 
        \DWACT_ADD_CI_0_g_array_0_1[0]\);
    
    un1_InitCnt_I_53 : XOR2
      port map(A => \InitCnt[2]_net_1\, B => \ClkEn\, Y => 
        \DWACT_ADD_CI_0_partial_sum[2]\);
    
    \InitCnt_RNO[5]\ : NOR2A
      port map(A => I_63, B => N_180, Y => \InitCnt_RNO[5]_net_1\);
    
    \DivCnt_RNIQ5QA[6]\ : NOR2B
      port map(A => \DivCnt[6]_net_1\, B => PAT_En, Y => 
        ClkEn_4_0_a4_0);
    
    un1_InitCnt_I_11 : AND2
      port map(A => \InitCnt[4]_net_1\, B => \ClkEn_0\, Y => 
        \DWACT_ADD_CI_0_g_array_0_4[0]\);
    
    \DivCnt[2]\ : DFN1C0
      port map(D => N_8, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \DivCnt[2]_net_1\);
    
    un1_InitCnt_I_90 : AO1
      port map(A => \DWACT_ADD_CI_0_pog_array_0_3[0]\, B => 
        \DWACT_ADD_CI_0_g_array_2[0]\, C => 
        \DWACT_ADD_CI_0_g_array_0_4[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_12_1[0]\);
    
    un1_InitCnt_I_40 : XOR2
      port map(A => \InitCnt[17]_net_1\, B => \ClkEn_1\, Y => 
        \DWACT_ADD_CI_0_partial_sum[17]\);
    
    un1_InitCnt_I_6 : AND2
      port map(A => \InitCnt[6]_net_1\, B => \ClkEn\, Y => 
        \DWACT_ADD_CI_0_g_array_0_6[0]\);
    
    \InitCnt_RNI2M3Q[14]\ : NOR3A
      port map(A => un27_clken_0_a2_0_6, B => \InitCnt[15]_net_1\, 
        C => \InitCnt[14]_net_1\, Y => un27_clken_0_a2_0_9);
    
    un1_InitCnt_I_99 : AO1
      port map(A => \DWACT_ADD_CI_0_pog_array_1_1[0]\, B => 
        \DWACT_ADD_CI_0_g_array_2[0]\, C => 
        \DWACT_ADD_CI_0_g_array_1_2[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_11[0]\);
    
    un1_InitCnt_I_49 : XOR2
      port map(A => \InitCnt[8]_net_1\, B => \ClkEn\, Y => 
        \DWACT_ADD_CI_0_partial_sum[8]\);
    
    un1_InitCnt_I_97 : AO1
      port map(A => \DWACT_ADD_CI_0_pog_array_0_9[0]\, B => 
        \DWACT_ADD_CI_0_g_array_11_1[0]\, C => 
        \DWACT_ADD_CI_0_g_array_0_10[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_12_4[0]\);
    
    un1_InitCnt_I_47 : XOR2
      port map(A => \InitCnt[7]_net_1\, B => \ClkEn\, Y => 
        \DWACT_ADD_CI_0_partial_sum[7]\);
    
    un1_InitCnt_I_20 : AND2
      port map(A => \InitCnt[11]_net_1\, B => \ClkEn_0\, Y => 
        \DWACT_ADD_CI_0_g_array_0_11[0]\);
    
    un1_InitCnt_I_94 : AO1
      port map(A => \DWACT_ADD_CI_0_pog_array_0_7[0]\, B => 
        \DWACT_ADD_CI_0_g_array_3[0]\, C => 
        \DWACT_ADD_CI_0_g_array_0_8[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_12_3[0]\);
    
    un1_InitCnt_I_44 : XOR2
      port map(A => \InitCnt[0]_net_1\, B => \ClkEn\, Y => 
        \DWACT_ADD_CI_0_partial_sum[0]\);
    
    \InitCnt[16]\ : DFN1C0
      port map(D => \InitCnt_RNO[16]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \InitCnt[16]_net_1\);
    
    un1_InitCnt_I_103 : AO1
      port map(A => \DWACT_ADD_CI_0_pog_array_0_15[0]\, B => 
        \DWACT_ADD_CI_0_g_array_4[0]\, C => 
        \DWACT_ADD_CI_0_g_array_0_16[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_12_7[0]\);
    
    un1_InitCnt_I_29 : XOR2
      port map(A => \InitCnt[3]_net_1\, B => \ClkEn_1\, Y => 
        \DWACT_ADD_CI_0_pog_array_0_2[0]\);
    
    \InitCnt_RNO[1]\ : NOR2A
      port map(A => I_62, B => N_180, Y => \InitCnt_RNO[1]_net_1\);
    
    un1_InitCnt_I_27 : XOR2
      port map(A => \InitCnt[10]_net_1\, B => \ClkEn_1\, Y => 
        \DWACT_ADD_CI_0_pog_array_0_9[0]\);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    \DivCnt_RNO[3]\ : XA1
      port map(A => \DivCnt[3]_net_1\, B => N_18, C => PAT_En, Y
         => N_10);
    
    \InitCnt_RNI5B2C[12]\ : NOR2
      port map(A => \InitCnt[12]_net_1\, B => \InitCnt[13]_net_1\, 
        Y => un27_clken_0_a2_0_4);
    
    \DivCnt_RNO_0[6]\ : NOR2B
      port map(A => N_20, B => \DivCnt[5]_net_1\, Y => N_171);
    
    un1_InitCnt_I_80 : AO1
      port map(A => \DWACT_ADD_CI_0_pog_array_0_10[0]\, B => 
        \DWACT_ADD_CI_0_g_array_0_10[0]\, C => 
        \DWACT_ADD_CI_0_g_array_0_11[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_1_5[0]\);
    
    un1_InitCnt_I_24 : XOR2
      port map(A => \InitCnt[6]_net_1\, B => \ClkEn_1\, Y => 
        \DWACT_ADD_CI_0_pog_array_0_5[0]\);
    
    mem_HL_RNO_0 : AO1D
      port map(A => un27_clken_0_a2_0, B => N_47, C => N_80, Y
         => un27_clken_0_o2_0);
    
    un1_InitCnt_I_30 : XOR2
      port map(A => \InitCnt[12]_net_1\, B => \ClkEn_1\, Y => 
        \DWACT_ADD_CI_0_pog_array_0_11[0]\);
    
    \InitCnt_RNI6LQ7_0[1]\ : NOR3
      port map(A => \InitCnt[1]_net_1\, B => N_47, C => 
        \InitCnt[4]_net_1\, Y => un1_pat_en_1_0_a2_0);
    
    un1_InitCnt_I_89 : AO1
      port map(A => \DWACT_ADD_CI_0_pog_array_1_4[0]\, B => 
        \DWACT_ADD_CI_0_g_array_1_4[0]\, C => 
        \DWACT_ADD_CI_0_g_array_1_5[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_2_2[0]\);
    
    \InitCnt_RNO[13]\ : NOR2A
      port map(A => I_58, B => N_180, Y => 
        \InitCnt_RNO[13]_net_1\);
    
    \DivCnt_RNI5VHP[3]\ : NOR3A
      port map(A => DivCnt_n1_0_i_a2_2, B => \DivCnt[4]_net_1\, C
         => \DivCnt[3]_net_1\, Y => N_41);
    
    un1_InitCnt_I_87 : AO1
      port map(A => \DWACT_ADD_CI_0_pog_array_0_13[0]\, B => 
        \DWACT_ADD_CI_0_g_array_11_2[0]\, C => 
        \DWACT_ADD_CI_0_g_array_0_14[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_12_6[0]\);
    
    un1_InitCnt_I_70 : XOR2
      port map(A => \DWACT_ADD_CI_0_partial_sum[9]\, B => 
        \DWACT_ADD_CI_0_g_array_12_3[0]\, Y => I_70);
    
    un1_InitCnt_I_95 : AO1
      port map(A => \DWACT_ADD_CI_0_pog_array_3[0]\, B => 
        \DWACT_ADD_CI_0_g_array_3[0]\, C => 
        \DWACT_ADD_CI_0_g_array_3_1[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_4[0]\);
    
    un1_InitCnt_I_39 : XOR2
      port map(A => \InitCnt[11]_net_1\, B => \ClkEn_1\, Y => 
        \DWACT_ADD_CI_0_partial_sum[11]\);
    
    un1_InitCnt_I_45 : XOR2
      port map(A => \InitCnt[12]_net_1\, B => \ClkEn\, Y => 
        \DWACT_ADD_CI_0_partial_sum[12]\);
    
    un1_InitCnt_I_96 : AO1
      port map(A => \DWACT_ADD_CI_0_pog_array_1[0]\, B => 
        \DWACT_ADD_CI_0_g_array_1[0]\, C => 
        \DWACT_ADD_CI_0_g_array_1_1[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_2[0]\);
    
    un1_InitCnt_I_37 : XOR2
      port map(A => \InitCnt[8]_net_1\, B => \ClkEn_1\, Y => 
        \DWACT_ADD_CI_0_pog_array_0_7[0]\);
    
    un1_InitCnt_I_46 : XOR2
      port map(A => \InitCnt[1]_net_1\, B => \ClkEn\, Y => 
        \DWACT_ADD_CI_0_partial_sum[1]\);
    
    \InitCnt_RNO[8]\ : NOR2A
      port map(A => I_69, B => N_180, Y => \InitCnt_RNO[8]_net_1\);
    
    \InitCnt_RNO[17]\ : NOR2A
      port map(A => I_74, B => N_180, Y => 
        \InitCnt_RNO[17]_net_1\);
    
    un1_InitCnt_I_84 : AO1
      port map(A => \DWACT_ADD_CI_0_pog_array_0_12[0]\, B => 
        \DWACT_ADD_CI_0_g_array_0_12[0]\, C => 
        \DWACT_ADD_CI_0_g_array_0_13[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_1_6[0]\);
    
    un1_InitCnt_I_42 : XOR2
      port map(A => \InitCnt[5]_net_1\, B => \ClkEn\, Y => 
        \DWACT_ADD_CI_0_partial_sum[5]\);
    
    un1_InitCnt_I_106 : AND2
      port map(A => \DWACT_ADD_CI_0_pog_array_0_7[0]\, B => 
        \DWACT_ADD_CI_0_pog_array_0_8[0]\, Y => 
        \DWACT_ADD_CI_0_pog_array_1_3[0]\);
    
    un1_InitCnt_I_105 : AND2
      port map(A => \DWACT_ADD_CI_0_pog_array_0_1[0]\, B => 
        \DWACT_ADD_CI_0_pog_array_0_2[0]\, Y => 
        \DWACT_ADD_CI_0_pog_array_1[0]\);
    
    un1_InitCnt_I_79 : AO1
      port map(A => \DWACT_ADD_CI_0_pog_array_1_6[0]\, B => 
        \DWACT_ADD_CI_0_g_array_1_6[0]\, C => 
        \DWACT_ADD_CI_0_g_array_1_7[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_2_3[0]\);
    
    un1_InitCnt_I_77 : AO1
      port map(A => \DWACT_ADD_CI_0_pog_array_0_2[0]\, B => 
        \DWACT_ADD_CI_0_g_array_0_2[0]\, C => 
        \DWACT_ADD_CI_0_g_array_0_3[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_1_1[0]\);
    
    un1_InitCnt_I_34 : XOR2
      port map(A => \InitCnt[9]_net_1\, B => \ClkEn_1\, Y => 
        \DWACT_ADD_CI_0_pog_array_0_8[0]\);
    
    \InitCnt[7]\ : DFN1C0
      port map(D => N_44, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \InitCnt[7]_net_1\);
    
    \InitCnt[3]\ : DFN1C0
      port map(D => \InitCnt_RNO[3]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \InitCnt[3]_net_1\);
    
    \DivCnt_RNIT57A[1]\ : NOR2B
      port map(A => \DivCnt[1]_net_1\, B => \DivCnt[0]_net_1\, Y
         => N_17);
    
    \DivCnt_RNO[0]\ : NOR2A
      port map(A => PAT_En, B => \DivCnt[0]_net_1\, Y => 
        DivCnt_n0);
    
    un1_InitCnt_I_68 : XOR2
      port map(A => \DWACT_ADD_CI_0_partial_sum[2]\, B => 
        \DWACT_ADD_CI_0_g_array_1[0]\, Y => I_68);
    
    un1_InitCnt_I_25 : XOR2
      port map(A => \InitCnt[13]_net_1\, B => \ClkEn_1\, Y => 
        \DWACT_ADD_CI_0_pog_array_0_12[0]\);
    
    \InitCnt_RNO[6]\ : NOR2A
      port map(A => I_65, B => N_180, Y => \InitCnt_RNO[6]_net_1\);
    
    un1_InitCnt_I_74 : XOR2
      port map(A => \DWACT_ADD_CI_0_partial_sum[17]\, B => 
        \DWACT_ADD_CI_0_g_array_12_7[0]\, Y => I_74);
    
    un1_InitCnt_I_26 : XOR2
      port map(A => \InitCnt[1]_net_1\, B => \ClkEn_1\, Y => 
        \DWACT_ADD_CI_0_pog_array_0[0]\);
    
    un1_InitCnt_I_101 : AO1
      port map(A => \DWACT_ADD_CI_0_pog_array_0_1[0]\, B => 
        \DWACT_ADD_CI_0_g_array_1[0]\, C => 
        \DWACT_ADD_CI_0_g_array_0_2[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_12[0]\);
    
    un1_InitCnt_I_22 : XOR2
      port map(A => \InitCnt[15]_net_1\, B => \ClkEn_1\, Y => 
        \DWACT_ADD_CI_0_pog_array_0_14[0]\);
    
    un1_InitCnt_I_61 : XOR2
      port map(A => \DWACT_ADD_CI_0_partial_sum[4]\, B => 
        \DWACT_ADD_CI_0_g_array_2[0]\, Y => I_61);
    
    \InitCnt_RNIQ5T7[6]\ : NOR3A
      port map(A => un27_clken_0_a2_0_2, B => \InitCnt[7]_net_1\, 
        C => \InitCnt[6]_net_1\, Y => un27_clken_0_a2_0_7);
    
    \DivCnt_RNO[6]\ : XA1B
      port map(A => \DivCnt[6]_net_1\, B => N_171, C => 
        DivCnt_n6_0_i_0, Y => N_16);
    
    un1_InitCnt_I_10 : AND2
      port map(A => \InitCnt[10]_net_1\, B => \ClkEn_0\, Y => 
        \DWACT_ADD_CI_0_g_array_0_10[0]\);
    
    un1_InitCnt_I_85 : AO1
      port map(A => \DWACT_ADD_CI_0_pog_array_0_6[0]\, B => 
        \DWACT_ADD_CI_0_g_array_0_6[0]\, C => 
        \DWACT_ADD_CI_0_g_array_0_7[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_1_3[0]\);
    
    \DivCnt_RNO[5]\ : XA1
      port map(A => \DivCnt[5]_net_1\, B => N_20, C => PAT_En, Y
         => N_14);
    
    un1_InitCnt_I_5 : AND2
      port map(A => \InitCnt[12]_net_1\, B => \ClkEn\, Y => 
        \DWACT_ADD_CI_0_g_array_0_12[0]\);
    
    un1_InitCnt_I_82 : AO1
      port map(A => \DWACT_ADD_CI_0_pog_array_1_3[0]\, B => 
        \DWACT_ADD_CI_0_g_array_3[0]\, C => 
        \DWACT_ADD_CI_0_g_array_1_4[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_11_1[0]\);
    
    un1_InitCnt_I_35 : XOR2
      port map(A => \InitCnt[7]_net_1\, B => \ClkEn_1\, Y => 
        \DWACT_ADD_CI_0_pog_array_0_6[0]\);
    
    un1_InitCnt_I_36 : XOR2
      port map(A => \InitCnt[16]_net_1\, B => \ClkEn_1\, Y => 
        \DWACT_ADD_CI_0_pog_array_0_15[0]\);
    
    un1_InitCnt_I_32 : XOR2
      port map(A => \InitCnt[2]_net_1\, B => \ClkEn_1\, Y => 
        \DWACT_ADD_CI_0_pog_array_0_1[0]\);
    
    un1_InitCnt_I_19 : AND2
      port map(A => \InitCnt[8]_net_1\, B => \ClkEn_0\, Y => 
        \DWACT_ADD_CI_0_g_array_0_8[0]\);
    
    un1_InitCnt_I_17 : AND2
      port map(A => \InitCnt[7]_net_1\, B => \ClkEn_0\, Y => 
        \DWACT_ADD_CI_0_g_array_0_7[0]\);
    
    un1_InitCnt_I_75 : AO1
      port map(A => \DWACT_ADD_CI_0_pog_array_0[0]\, B => 
        \DWACT_ADD_CI_0_TMP[0]\, C => 
        \DWACT_ADD_CI_0_g_array_0_1[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_1[0]\);
    
    \InitCnt_RNINGPB[0]\ : OR3B
      port map(A => PAT_En, B => \ClkEn_0\, C => 
        \InitCnt[0]_net_1\, Y => \InitCnt_5_i_a3_1[0]\);
    
    \InitCnt_RNO[15]\ : NOR2A
      port map(A => I_66, B => N_180, Y => 
        \InitCnt_RNO[15]_net_1\);
    
    un1_InitCnt_I_76 : AO1
      port map(A => \DWACT_ADD_CI_0_pog_array_0_8[0]\, B => 
        \DWACT_ADD_CI_0_g_array_0_8[0]\, C => 
        \DWACT_ADD_CI_0_g_array_0_9[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_1_4[0]\);
    
    reset_RNO : AO1B
      port map(A => un1_pat_en_1_0_a2_0, B => N_94, C => PAT_En, 
        Y => un1_pat_en_1);
    
    un1_InitCnt_I_72 : XOR2
      port map(A => \DWACT_ADD_CI_0_partial_sum[3]\, B => 
        \DWACT_ADD_CI_0_g_array_12[0]\, Y => I_72);
    
    mem_HL_RNO_2 : NOR3B
      port map(A => \InitCnt[0]_net_1\, B => \InitCnt[1]_net_1\, 
        C => \InitCnt[4]_net_1\, Y => N_80);
    
    un1_InitCnt_I_14 : AND2
      port map(A => \InitCnt[14]_net_1\, B => \ClkEn_0\, Y => 
        \DWACT_ADD_CI_0_g_array_0_14[0]\);
    
    ClkEn_0 : DFN1C0
      port map(D => ClkEn_4, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \ClkEn_0\);
    
    precharge : DFN1E1P0
      port map(D => un39_clken, CLK => PLL_Test1_0_Sys_66M_Clk, 
        PRE => PLL_Test1_0_SysRst_O, E => \ClkEn_0\, Q => 
        precharge_c);
    
    \InitCnt_RNO[7]\ : OA1A
      port map(A => PAT_En, B => I_67, C => N_73, Y => N_44);
    
    \InitCnt_RNO[9]\ : NOR2A
      port map(A => I_70, B => N_180, Y => \InitCnt_RNO[9]_net_1\);
    
    \InitCnt_RNO[14]\ : NOR2A
      port map(A => I_64, B => N_180, Y => 
        \InitCnt_RNO[14]_net_1\);
    
    \InitCnt_RNO[3]\ : OA1A
      port map(A => PAT_En, B => I_72, C => N_73, Y => 
        \InitCnt_RNO[3]_net_1\);
    
    \InitCnt_RNIPA1E[17]\ : NOR3
      port map(A => \InitCnt[5]_net_1\, B => \InitCnt[17]_net_1\, 
        C => \InitCnt[16]_net_1\, Y => un27_clken_0_a2_0_6);
    
    \InitCnt[12]\ : DFN1C0
      port map(D => \InitCnt_RNO[12]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \InitCnt[12]_net_1\);
    
    un1_InitCnt_I_93 : AO1
      port map(A => \DWACT_ADD_CI_0_pog_array_0_5[0]\, B => 
        \DWACT_ADD_CI_0_g_array_11[0]\, C => 
        \DWACT_ADD_CI_0_g_array_0_6[0]\, Y => 
        \DWACT_ADD_CI_0_g_array_12_2[0]\);
    
    un1_InitCnt_I_43 : XOR2
      port map(A => \InitCnt[13]_net_1\, B => \ClkEn\, Y => 
        \DWACT_ADD_CI_0_partial_sum[13]\);
    
    \InitCnt[14]\ : DFN1C0
      port map(D => \InitCnt_RNO[14]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \InitCnt[14]_net_1\);
    
    mem_HL_RNO_1 : OR2A
      port map(A => \InitCnt[4]_net_1\, B => \InitCnt[0]_net_1\, 
        Y => un27_clken_0_a2_0);
    
    \InitCnt_RNI95382[0]\ : OR3B
      port map(A => N_94, B => un1_pat_en_1_0_a2_0, C => 
        un1_initcnt14_i_a3_0, Y => N_69);
    
    un1_InitCnt_I_15 : AND2
      port map(A => \InitCnt[15]_net_1\, B => \ClkEn_0\, Y => 
        \DWACT_ADD_CI_0_g_array_0_15[0]\);
    
    un1_InitCnt_I_16 : AND2
      port map(A => \InitCnt[13]_net_1\, B => \ClkEn_0\, Y => 
        \DWACT_ADD_CI_0_g_array_0_13[0]\);
    
    \InitCnt_RNI6M4O[10]\ : NOR3A
      port map(A => un27_clken_0_a2_0_4, B => \InitCnt[11]_net_1\, 
        C => \InitCnt[10]_net_1\, Y => un27_clken_0_a2_0_8);
    
    un1_InitCnt_I_12 : AND2
      port map(A => \InitCnt[2]_net_1\, B => \ClkEn_0\, Y => 
        \DWACT_ADD_CI_0_g_array_0_2[0]\);
    
    un1_InitCnt_I_23 : XOR2
      port map(A => \InitCnt[4]_net_1\, B => \ClkEn_1\, Y => 
        \DWACT_ADD_CI_0_pog_array_0_3[0]\);
    
    \DivCnt[3]\ : DFN1C0
      port map(D => N_10, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \DivCnt[3]_net_1\);
    
    \DivCnt_RNO_0[1]\ : XAI1
      port map(A => \DivCnt[0]_net_1\, B => \DivCnt[1]_net_1\, C
         => PAT_En, Y => DivCnt_n1_0_i_1);
    
    \InitCnt[9]\ : DFN1C0
      port map(D => \InitCnt_RNO[9]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \InitCnt[9]_net_1\);
    
    mem_HL : DFN1E1P0
      port map(D => un27_clken, CLK => PLL_Test1_0_Sys_66M_Clk, 
        PRE => PLL_Test1_0_SysRst_O, E => \ClkEn_0\, Q => 
        mem_HL_c);
    
    un1_InitCnt_I_58 : XOR2
      port map(A => \DWACT_ADD_CI_0_partial_sum[13]\, B => 
        \DWACT_ADD_CI_0_g_array_12_5[0]\, Y => I_58);
    
    \DivCnt[6]\ : DFN1C0
      port map(D => N_16, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \DivCnt[6]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3;
use proasic3.all;

entity CMOS_DrvX is

    port( CMOS_reset_c             : out   std_logic;
          CMOS_sample_c            : out   std_logic;
          precharge_c              : out   std_logic;
          mem_HL_c                 : out   std_logic;
          spi_load_c               : out   std_logic;
          spi_data_c               : out   std_logic;
          spi_clock_c              : out   std_logic;
          CMOS_DrvX_VCC            : in    std_logic;
          PLL_Test1_0_ADC_66M_Clk  : in    std_logic;
          DRY_c_c                  : out   std_logic;
          CMOS_DrvX_0_AdcEn        : out   std_logic;
          Sync_Y_c                 : out   std_logic;
          Clock_Y_c                : out   std_logic;
          NoRowSel_c               : out   std_logic;
          Pre_co_c                 : out   std_logic;
          Sh_co_c                  : out   std_logic;
          Sync_X_c                 : out   std_logic;
          Clock_X_c                : out   std_logic;
          CMOS_DrvX_0_LVDSen_3     : out   std_logic;
          PLL_Test1_0_Sys_66M_Clk  : in    std_logic;
          PLL_Test1_0_SysRst_O     : in    std_logic;
          CMOS_DrvX_0_LVDSen_2     : out   std_logic;
          CMOS_DrvX_0_LVDSen_1     : out   std_logic;
          CMOS_DrvX_0_LVDSen_0     : out   std_logic;
          CMOS_DrvX_0_SDramEn_5    : out   std_logic;
          CMOS_DrvX_0_SDramEn_4    : out   std_logic;
          CMOS_DrvX_0_SDramEn_3    : out   std_logic;
          CMOS_DrvX_0_SDramEn_2    : out   std_logic;
          CMOS_DrvX_0_SDramEn_1    : out   std_logic;
          CMOS_DrvX_0_SDramEn_0    : out   std_logic;
          Sdram_cmd_0_SDoneFrameOk : in    std_logic;
          FrameMk_0_LVDS_ok        : in    std_logic;
          CMOS_DrvX_0_LVDSen       : out   std_logic;
          CMOS_DrvX_0_SDramEn      : out   std_logic;
          CMOS_DrvX_GND            : in    std_logic
        );

end CMOS_DrvX;

architecture DEF_ARCH of CMOS_DrvX is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component Y_X_Addressing
    port( Clock_X_c               : out   std_logic;
          Sync_X_c                : out   std_logic;
          Sh_co_c                 : out   std_logic;
          Pre_co_c                : out   std_logic;
          NoRowSel_c              : out   std_logic;
          Clock_Y_c               : out   std_logic;
          Sync_Y_c                : out   std_logic;
          CMOS_DrvX_0_AdcEn       : out   std_logic;
          ImageOrQl               : in    std_logic := 'U';
          DRY_c_c                 : out   std_logic;
          PLL_Test1_0_ADC_66M_Clk : in    std_logic := 'U';
          Y_X_Addressing_GND      : in    std_logic := 'U';
          Y_X_Addressing_VCC      : in    std_logic := 'U';
          Y_X_WaveEn_i            : in    std_logic := 'U';
          Y_X_WaveOk              : out   std_logic;
          Y_X_WaveEn              : in    std_logic := 'U';
          PLL_Test1_0_SysRst_O    : in    std_logic := 'U';
          PLL_Test1_0_Sys_66M_Clk : in    std_logic := 'U'
        );
  end component;

  component CMOS_Ctl
    port( CMOS_Ctl_GND             : in    std_logic := 'U';
          CMOS_DrvX_0_SDramEn      : out   std_logic;
          ImageOrQl                : out   std_logic;
          SPI_En                   : out   std_logic;
          PAT_En                   : out   std_logic;
          CMOS_DrvX_0_LVDSen       : out   std_logic;
          FrameMk_0_LVDS_ok        : in    std_logic := 'U';
          Sdram_cmd_0_SDoneFrameOk : in    std_logic := 'U';
          Y_X_WaveOk               : in    std_logic := 'U';
          PAT_Ok                   : in    std_logic := 'U';
          SPI_Ok                   : in    std_logic := 'U';
          SPI_En_i                 : out   std_logic;
          Y_X_WaveEn               : out   std_logic;
          Y_X_WaveEn_i             : out   std_logic;
          SPI_En_0                 : out   std_logic;
          CMOS_DrvX_0_SDramEn_0    : out   std_logic;
          CMOS_DrvX_0_SDramEn_1    : out   std_logic;
          CMOS_DrvX_0_SDramEn_2    : out   std_logic;
          CMOS_DrvX_0_SDramEn_3    : out   std_logic;
          CMOS_DrvX_0_SDramEn_4    : out   std_logic;
          CMOS_DrvX_0_SDramEn_5    : out   std_logic;
          CMOS_DrvX_0_LVDSen_0     : out   std_logic;
          CMOS_DrvX_0_LVDSen_1     : out   std_logic;
          CMOS_DrvX_0_LVDSen_2     : out   std_logic;
          PLL_Test1_0_SysRst_O     : in    std_logic := 'U';
          PLL_Test1_0_Sys_66M_Clk  : in    std_logic := 'U';
          CMOS_DrvX_0_LVDSen_3     : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component SPI_Set
    port( SPI_En_i                : in    std_logic := 'U';
          spi_clock_c             : out   std_logic;
          spi_data_c              : out   std_logic;
          spi_load_c              : out   std_logic;
          SPI_Ok                  : out   std_logic;
          PLL_Test1_0_SysRst_O    : in    std_logic := 'U';
          PLL_Test1_0_Sys_66M_Clk : in    std_logic := 'U';
          SPI_En                  : in    std_logic := 'U';
          SPI_En_0                : in    std_logic := 'U'
        );
  end component;

  component PixelArrayTiming
    port( PAT_Ok                  : out   std_logic;
          mem_HL_c                : out   std_logic;
          precharge_c             : out   std_logic;
          CMOS_sample_c           : out   std_logic;
          CMOS_reset_c            : out   std_logic;
          PAT_En                  : in    std_logic := 'U';
          PLL_Test1_0_SysRst_O    : in    std_logic := 'U';
          PLL_Test1_0_Sys_66M_Clk : in    std_logic := 'U'
        );
  end component;

    signal ImageOrQl, SPI_En, PAT_En, Y_X_WaveOk, PAT_Ok, SPI_Ok, 
        SPI_En_i, Y_X_WaveEn, Y_X_WaveEn_i, SPI_En_0, \GND\, 
        \VCC\, GND_0, VCC_0 : std_logic;

    for all : Y_X_Addressing
	Use entity work.Y_X_Addressing(DEF_ARCH);
    for all : CMOS_Ctl
	Use entity work.CMOS_Ctl(DEF_ARCH);
    for all : SPI_Set
	Use entity work.SPI_Set(DEF_ARCH);
    for all : PixelArrayTiming
	Use entity work.PixelArrayTiming(DEF_ARCH);
begin 


    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    Module_Y_X_Addressing : Y_X_Addressing
      port map(Clock_X_c => Clock_X_c, Sync_X_c => Sync_X_c, 
        Sh_co_c => Sh_co_c, Pre_co_c => Pre_co_c, NoRowSel_c => 
        NoRowSel_c, Clock_Y_c => Clock_Y_c, Sync_Y_c => Sync_Y_c, 
        CMOS_DrvX_0_AdcEn => CMOS_DrvX_0_AdcEn, ImageOrQl => 
        ImageOrQl, DRY_c_c => DRY_c_c, PLL_Test1_0_ADC_66M_Clk
         => PLL_Test1_0_ADC_66M_Clk, Y_X_Addressing_GND => 
        CMOS_DrvX_GND, Y_X_Addressing_VCC => CMOS_DrvX_VCC, 
        Y_X_WaveEn_i => Y_X_WaveEn_i, Y_X_WaveOk => Y_X_WaveOk, 
        Y_X_WaveEn => Y_X_WaveEn, PLL_Test1_0_SysRst_O => 
        PLL_Test1_0_SysRst_O, PLL_Test1_0_Sys_66M_Clk => 
        PLL_Test1_0_Sys_66M_Clk);
    
    Module_CMOS_Ctl : CMOS_Ctl
      port map(CMOS_Ctl_GND => CMOS_DrvX_GND, CMOS_DrvX_0_SDramEn
         => CMOS_DrvX_0_SDramEn, ImageOrQl => ImageOrQl, SPI_En
         => SPI_En, PAT_En => PAT_En, CMOS_DrvX_0_LVDSen => 
        CMOS_DrvX_0_LVDSen, FrameMk_0_LVDS_ok => 
        FrameMk_0_LVDS_ok, Sdram_cmd_0_SDoneFrameOk => 
        Sdram_cmd_0_SDoneFrameOk, Y_X_WaveOk => Y_X_WaveOk, 
        PAT_Ok => PAT_Ok, SPI_Ok => SPI_Ok, SPI_En_i => SPI_En_i, 
        Y_X_WaveEn => Y_X_WaveEn, Y_X_WaveEn_i => Y_X_WaveEn_i, 
        SPI_En_0 => SPI_En_0, CMOS_DrvX_0_SDramEn_0 => 
        CMOS_DrvX_0_SDramEn_0, CMOS_DrvX_0_SDramEn_1 => 
        CMOS_DrvX_0_SDramEn_1, CMOS_DrvX_0_SDramEn_2 => 
        CMOS_DrvX_0_SDramEn_2, CMOS_DrvX_0_SDramEn_3 => 
        CMOS_DrvX_0_SDramEn_3, CMOS_DrvX_0_SDramEn_4 => 
        CMOS_DrvX_0_SDramEn_4, CMOS_DrvX_0_SDramEn_5 => 
        CMOS_DrvX_0_SDramEn_5, CMOS_DrvX_0_LVDSen_0 => 
        CMOS_DrvX_0_LVDSen_0, CMOS_DrvX_0_LVDSen_1 => 
        CMOS_DrvX_0_LVDSen_1, CMOS_DrvX_0_LVDSen_2 => 
        CMOS_DrvX_0_LVDSen_2, PLL_Test1_0_SysRst_O => 
        PLL_Test1_0_SysRst_O, PLL_Test1_0_Sys_66M_Clk => 
        PLL_Test1_0_Sys_66M_Clk, CMOS_DrvX_0_LVDSen_3 => 
        CMOS_DrvX_0_LVDSen_3);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    Module_SPI_Set : SPI_Set
      port map(SPI_En_i => SPI_En_i, spi_clock_c => spi_clock_c, 
        spi_data_c => spi_data_c, spi_load_c => spi_load_c, 
        SPI_Ok => SPI_Ok, PLL_Test1_0_SysRst_O => 
        PLL_Test1_0_SysRst_O, PLL_Test1_0_Sys_66M_Clk => 
        PLL_Test1_0_Sys_66M_Clk, SPI_En => SPI_En, SPI_En_0 => 
        SPI_En_0);
    
    Module_PixelArrayTiming : PixelArrayTiming
      port map(PAT_Ok => PAT_Ok, mem_HL_c => mem_HL_c, 
        precharge_c => precharge_c, CMOS_sample_c => 
        CMOS_sample_c, CMOS_reset_c => CMOS_reset_c, PAT_En => 
        PAT_En, PLL_Test1_0_SysRst_O => PLL_Test1_0_SysRst_O, 
        PLL_Test1_0_Sys_66M_Clk => PLL_Test1_0_Sys_66M_Clk);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3;
use proasic3.all;

entity My_adder0 is

    port( intData2acc_RNICNV9                         : in    std_logic_vector(46 to 46);
          intData2acc_RNIBNV9                         : in    std_logic_vector(45 to 45);
          intData2acc_RNI9RV9                         : in    std_logic_vector(51 to 51);
          intData2acc_RNI6JV9                         : in    std_logic_vector(36 to 36);
          intData2acc_RNI7JV9                         : in    std_logic_vector(37 to 37);
          intData2acc_RNI6NV9                         : in    std_logic_vector(40 to 40);
          intData2acc_RNIENV9                         : in    std_logic_vector(48 to 48);
          intData2acc_RNI8RV9                         : in    std_logic_vector(50 to 50);
          intData2acc_RNIBJV9                         : in    std_logic_vector(38 to 38);
          intData2acc_RNICJV9                         : in    std_logic_vector(39 to 39);
          intData2acc_RNIFNV9                         : in    std_logic_vector(49 to 49);
          intData2acc_RNI8NV9                         : in    std_logic_vector(42 to 42);
          intData2acc_RNI9NV9                         : in    std_logic_vector(43 to 43);
          intData2acc_RNIDNV9                         : in    std_logic_vector(47 to 47);
          intData2acc_RNI7NV9                         : in    std_logic_vector(41 to 41);
          intData2acc_RNIANV9                         : in    std_logic_vector(44 to 44);
          intData2acc_RNIBRV9                         : in    std_logic_vector(53 downto 52);
          \Z\\My_adder0_2_Sum_[15]\\\                 : out   std_logic;
          \Z\\My_adder0_2_Sum_[12]\\\                 : out   std_logic;
          \Z\\My_adder0_2_Sum_[6]\\\                  : out   std_logic;
          \Z\\My_adder0_2_Sum_[10]\\\                 : out   std_logic;
          \Z\\My_adder0_2_Sum_[9]\\\                  : out   std_logic;
          \Z\\My_adder0_2_Sum_[7]\\\                  : out   std_logic;
          \Z\\My_adder0_2_Sum_[11]\\\                 : out   std_logic;
          \Z\\My_adder0_2_Sum_[1]\\\                  : out   std_logic;
          \Z\\My_adder0_2_Sum_[3]\\\                  : out   std_logic;
          \Z\\My_adder0_2_Sum_[13]\\\                 : out   std_logic;
          \Z\\My_adder0_2_Sum_[0]\\\                  : out   std_logic;
          \Z\\My_adder0_2_Sum_[8]\\\                  : out   std_logic;
          \Z\\My_adder0_2_Sum_[14]\\\                 : out   std_logic;
          \Z\\adc_muxtmp_test_0_DataOut41to28_[29]\\\ : in    std_logic;
          \Z\\My_adder0_2_Sum_[2]\\\                  : out   std_logic;
          \Z\\My_adder0_2_Sum_[4]\\\                  : out   std_logic;
          \Z\\My_adder0_2_Sum_[5]\\\                  : out   std_logic;
          \Z\\My_adder0_2_Sum_[17]\\\                 : out   std_logic;
          My_adder0_GND                               : in    std_logic;
          \Z\\My_adder0_2_Sum_[16]\\\                 : out   std_logic
        );

end My_adder0;

architecture DEF_ARCH of My_adder0 is 

  component XOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MAJ3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component AND2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal Carry_15_net, Carry_8_net, Carry_7_net, Carry_5_net, 
        Carry_4_net, Carry_16_net, Carry_11_net, Carry_10_net, 
        Carry_6_net, Carry_13_net, Carry_12_net, Carry_3_net, 
        Carry_2_net, Carry_1_net, Carry_14_net, Carry_0_net, 
        Carry_9_net, \GND\, \VCC\, GND_0, VCC_0 : std_logic;

begin 


    XOR3_Sum_16_inst : XOR3
      port map(A => My_adder0_GND, B => intData2acc_RNIBRV9(52), 
        C => Carry_15_net, Y => \Z\\My_adder0_2_Sum_[16]\\\);
    
    MAJ3_Carry_8_inst : MAJ3
      port map(A => Carry_7_net, B => My_adder0_GND, C => 
        intData2acc_RNIANV9(44), Y => Carry_8_net);
    
    MAJ3_Carry_9_inst : MAJ3
      port map(A => Carry_8_net, B => My_adder0_GND, C => 
        intData2acc_RNIBNV9(45), Y => Carry_9_net);
    
    XOR3_Sum_5_inst : XOR3
      port map(A => My_adder0_GND, B => intData2acc_RNI7NV9(41), 
        C => Carry_4_net, Y => \Z\\My_adder0_2_Sum_[5]\\\);
    
    XOR3_Sum_2_inst : XOR3
      port map(A => My_adder0_GND, B => intData2acc_RNIBJV9(38), 
        C => Carry_1_net, Y => \Z\\My_adder0_2_Sum_[2]\\\);
    
    XOR3_Sum_4_inst : XOR3
      port map(A => My_adder0_GND, B => intData2acc_RNI6NV9(40), 
        C => Carry_3_net, Y => \Z\\My_adder0_2_Sum_[4]\\\);
    
    XOR3_Sum_11_inst : XOR3
      port map(A => My_adder0_GND, B => intData2acc_RNIDNV9(47), 
        C => Carry_10_net, Y => \Z\\My_adder0_2_Sum_[11]\\\);
    
    XOR3_Sum_12_inst : XOR3
      port map(A => My_adder0_GND, B => intData2acc_RNIENV9(48), 
        C => Carry_11_net, Y => \Z\\My_adder0_2_Sum_[12]\\\);
    
    MAJ3_Carry_5_inst : MAJ3
      port map(A => Carry_4_net, B => My_adder0_GND, C => 
        intData2acc_RNI7NV9(41), Y => Carry_5_net);
    
    MAJ3_Carry_2_inst : MAJ3
      port map(A => Carry_1_net, B => My_adder0_GND, C => 
        intData2acc_RNIBJV9(38), Y => Carry_2_net);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    MAJ3_Carry_1_inst : MAJ3
      port map(A => Carry_0_net, B => 
        \Z\\adc_muxtmp_test_0_DataOut41to28_[29]\\\, C => 
        intData2acc_RNI7JV9(37), Y => Carry_1_net);
    
    MAJ3_Carry_4_inst : MAJ3
      port map(A => Carry_3_net, B => My_adder0_GND, C => 
        intData2acc_RNI6NV9(40), Y => Carry_4_net);
    
    XOR3_Sum_13_inst : XOR3
      port map(A => My_adder0_GND, B => intData2acc_RNIFNV9(49), 
        C => Carry_12_net, Y => \Z\\My_adder0_2_Sum_[13]\\\);
    
    XOR3_Sum_1_inst : XOR3
      port map(A => \Z\\adc_muxtmp_test_0_DataOut41to28_[29]\\\, 
        B => intData2acc_RNI7JV9(37), C => Carry_0_net, Y => 
        \Z\\My_adder0_2_Sum_[1]\\\);
    
    MAJ3_Carry_12_inst : MAJ3
      port map(A => Carry_11_net, B => My_adder0_GND, C => 
        intData2acc_RNIENV9(48), Y => Carry_12_net);
    
    XOR3_Sum_17_inst : XOR3
      port map(A => My_adder0_GND, B => intData2acc_RNIBRV9(53), 
        C => Carry_16_net, Y => \Z\\My_adder0_2_Sum_[17]\\\);
    
    MAJ3_Carry_7_inst : MAJ3
      port map(A => Carry_6_net, B => My_adder0_GND, C => 
        intData2acc_RNI9NV9(43), Y => Carry_7_net);
    
    GND_i : GND
      port map(Y => \GND\);
    
    XOR3_Sum_6_inst : XOR3
      port map(A => My_adder0_GND, B => intData2acc_RNI8NV9(42), 
        C => Carry_5_net, Y => \Z\\My_adder0_2_Sum_[6]\\\);
    
    MAJ3_Carry_14_inst : MAJ3
      port map(A => Carry_13_net, B => My_adder0_GND, C => 
        intData2acc_RNI8RV9(50), Y => Carry_14_net);
    
    MAJ3_Carry_13_inst : MAJ3
      port map(A => Carry_12_net, B => My_adder0_GND, C => 
        intData2acc_RNIFNV9(49), Y => Carry_13_net);
    
    XOR3_Sum_3_inst : XOR3
      port map(A => My_adder0_GND, B => intData2acc_RNICJV9(39), 
        C => Carry_2_net, Y => \Z\\My_adder0_2_Sum_[3]\\\);
    
    XOR3_Sum_14_inst : XOR3
      port map(A => My_adder0_GND, B => intData2acc_RNI8RV9(50), 
        C => Carry_13_net, Y => \Z\\My_adder0_2_Sum_[14]\\\);
    
    XOR3_Sum_8_inst : XOR3
      port map(A => My_adder0_GND, B => intData2acc_RNIANV9(44), 
        C => Carry_7_net, Y => \Z\\My_adder0_2_Sum_[8]\\\);
    
    MAJ3_Carry_11_inst : MAJ3
      port map(A => Carry_10_net, B => My_adder0_GND, C => 
        intData2acc_RNIDNV9(47), Y => Carry_11_net);
    
    MAJ3_Carry_16_inst : MAJ3
      port map(A => Carry_15_net, B => My_adder0_GND, C => 
        intData2acc_RNIBRV9(52), Y => Carry_16_net);
    
    XOR3_Sum_7_inst : XOR3
      port map(A => My_adder0_GND, B => intData2acc_RNI9NV9(43), 
        C => Carry_6_net, Y => \Z\\My_adder0_2_Sum_[7]\\\);
    
    MAJ3_Carry_10_inst : MAJ3
      port map(A => Carry_9_net, B => My_adder0_GND, C => 
        intData2acc_RNICNV9(46), Y => Carry_10_net);
    
    MAJ3_Carry_3_inst : MAJ3
      port map(A => Carry_2_net, B => My_adder0_GND, C => 
        intData2acc_RNICJV9(39), Y => Carry_3_net);
    
    XOR3_Sum_15_inst : XOR3
      port map(A => My_adder0_GND, B => intData2acc_RNI9RV9(51), 
        C => Carry_14_net, Y => \Z\\My_adder0_2_Sum_[15]\\\);
    
    AND2_Carry_0_inst : AND2
      port map(A => My_adder0_GND, B => intData2acc_RNI6JV9(36), 
        Y => Carry_0_net);
    
    MAJ3_Carry_15_inst : MAJ3
      port map(A => Carry_14_net, B => My_adder0_GND, C => 
        intData2acc_RNI9RV9(51), Y => Carry_15_net);
    
    XOR3_Sum_9_inst : XOR3
      port map(A => My_adder0_GND, B => intData2acc_RNIBNV9(45), 
        C => Carry_8_net, Y => \Z\\My_adder0_2_Sum_[9]\\\);
    
    XOR2_Sum_0_inst : XOR2
      port map(A => My_adder0_GND, B => intData2acc_RNI6JV9(36), 
        Y => \Z\\My_adder0_2_Sum_[0]\\\);
    
    MAJ3_Carry_6_inst : MAJ3
      port map(A => Carry_5_net, B => My_adder0_GND, C => 
        intData2acc_RNI8NV9(42), Y => Carry_6_net);
    
    XOR3_Sum_10_inst : XOR3
      port map(A => My_adder0_GND, B => intData2acc_RNICNV9(46), 
        C => Carry_9_net, Y => \Z\\My_adder0_2_Sum_[10]\\\);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3;
use proasic3.all;

entity SDRAM_wr is

    port( \Z\\SDRAM_wr_0_wr_state_[2]\\\ : out   std_logic;
          \Z\\SDRAM_wr_0_wr_state_[1]\\\ : out   std_logic;
          \Z\\SDRAM_wr_0_wr_state_[0]\\\ : out   std_logic;
          Sdram_ctl_v2_0_SD_wrEn_i       : in    std_logic;
          PLL_Test1_0_SysRst_O           : in    std_logic;
          PLL_Test1_0_Sys_66M_Clk        : in    std_logic;
          SDRAM_wr_0_SD_WrOK             : out   std_logic;
          Sdram_cmd_0_wrrow_end          : in    std_logic;
          Sdram_ctl_v2_0_SD_wrEn         : in    std_logic
        );

end SDRAM_wr;

architecture DEF_ARCH of SDRAM_wr is 

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component XA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \wr_state_RNO[2]_net_1\, \pr_state[1]_net_1\, 
        \pr_state[0]_net_1\, \pr_state[2]_net_1\, 
        \wr_state_RNO[1]_net_1\, \pr_state[3]_net_1\, 
        \pr_state[4]_net_1\, \wr_state_RNO[0]_net_1\, 
        \pr_state[5]_net_1\, temp_n2, \temp[0]_net_1\, 
        \temp[1]_net_1\, N_25, N_90, \pr_state[6]_net_1\, N_73_i, 
        \temp[2]_net_1\, N_22, \pr_state_RNO_2[2]\, N_10, N_4, 
        temp_n0, N_39, N_69_i, N_67_i, \GND\, \VCC\, GND_0, VCC_0
         : std_logic;

begin 


    \wr_state[0]\ : DFN1C0
      port map(D => \wr_state_RNO[0]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \Z\\SDRAM_wr_0_wr_state_[0]\\\);
    
    \pr_state_RNO_0[5]\ : OR3B
      port map(A => \pr_state[6]_net_1\, B => 
        Sdram_ctl_v2_0_SD_wrEn, C => Sdram_cmd_0_wrrow_end, Y => 
        N_90);
    
    \wr_state_RNO[0]\ : OR3
      port map(A => \pr_state[1]_net_1\, B => \pr_state[5]_net_1\, 
        C => \pr_state[4]_net_1\, Y => \wr_state_RNO[0]_net_1\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    temp_n0_0_0_a3 : NOR2
      port map(A => \temp[0]_net_1\, B => N_25, Y => temp_n0);
    
    \pr_state_RNO[5]\ : AO1B
      port map(A => Sdram_ctl_v2_0_SD_wrEn, B => 
        \pr_state[0]_net_1\, C => N_90, Y => N_10);
    
    \wr_state_RNO[1]\ : OR3
      port map(A => \pr_state[0]_net_1\, B => \pr_state[3]_net_1\, 
        C => \pr_state[4]_net_1\, Y => \wr_state_RNO[1]_net_1\);
    
    \wr_state[1]\ : DFN1C0
      port map(D => \wr_state_RNO[1]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \Z\\SDRAM_wr_0_wr_state_[1]\\\);
    
    \pr_state[3]\ : DFN1C0
      port map(D => N_69_i, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \pr_state[3]_net_1\);
    
    wr_ok : DFN1C0
      port map(D => N_4, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => SDRAM_wr_0_SD_WrOK);
    
    \wr_state_RNO[2]\ : OR3
      port map(A => \pr_state[1]_net_1\, B => \pr_state[0]_net_1\, 
        C => \pr_state[2]_net_1\, Y => \wr_state_RNO[2]_net_1\);
    
    \temp[1]\ : DFN1C0
      port map(D => N_22, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \temp[1]_net_1\);
    
    wr_ok_RNO : NOR2B
      port map(A => \temp[2]_net_1\, B => \pr_state[2]_net_1\, Y
         => N_4);
    
    \pr_state[2]\ : DFN1C0
      port map(D => \pr_state_RNO_2[2]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \pr_state[2]_net_1\);
    
    \pr_state_RNO[0]\ : NOR2B
      port map(A => Sdram_ctl_v2_0_SD_wrEn, B => 
        \pr_state[1]_net_1\, Y => N_39);
    
    \temp[2]\ : DFN1C0
      port map(D => temp_n2, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \temp[2]_net_1\);
    
    temp_n1_0_i_o3 : OR2A
      port map(A => \pr_state[2]_net_1\, B => \temp[2]_net_1\, Y
         => N_25);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \pr_state_RNO[4]\ : NOR2B
      port map(A => Sdram_ctl_v2_0_SD_wrEn, B => 
        \pr_state[3]_net_1\, Y => N_67_i);
    
    \pr_state_RNO[1]\ : NOR3C
      port map(A => \pr_state[6]_net_1\, B => 
        Sdram_ctl_v2_0_SD_wrEn, C => Sdram_cmd_0_wrrow_end, Y => 
        N_73_i);
    
    temp_17_0_a3 : NOR3B
      port map(A => \temp[0]_net_1\, B => \temp[1]_net_1\, C => 
        N_25, Y => temp_n2);
    
    \pr_state[0]\ : DFN1C0
      port map(D => N_39, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \pr_state[0]_net_1\);
    
    \pr_state_RNO[2]\ : OA1
      port map(A => \pr_state[2]_net_1\, B => \pr_state[4]_net_1\, 
        C => Sdram_ctl_v2_0_SD_wrEn, Y => \pr_state_RNO_2[2]\);
    
    \temp[0]\ : DFN1C0
      port map(D => temp_n0, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \temp[0]_net_1\);
    
    \pr_state[4]\ : DFN1C0
      port map(D => N_67_i, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \pr_state[4]_net_1\);
    
    \pr_state[6]\ : DFN1P0
      port map(D => Sdram_ctl_v2_0_SD_wrEn_i, CLK => 
        PLL_Test1_0_Sys_66M_Clk, PRE => PLL_Test1_0_SysRst_O, Q
         => \pr_state[6]_net_1\);
    
    \pr_state[1]\ : DFN1C0
      port map(D => N_73_i, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \pr_state[1]_net_1\);
    
    \pr_state[5]\ : DFN1C0
      port map(D => N_10, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \pr_state[5]_net_1\);
    
    temp_n1_0_i : XA1B
      port map(A => \temp[0]_net_1\, B => \temp[1]_net_1\, C => 
        N_25, Y => N_22);
    
    \pr_state_RNO[3]\ : NOR2B
      port map(A => Sdram_ctl_v2_0_SD_wrEn, B => 
        \pr_state[5]_net_1\, Y => N_69_i);
    
    \wr_state[2]\ : DFN1C0
      port map(D => \wr_state_RNO[2]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \Z\\SDRAM_wr_0_wr_state_[2]\\\);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3;
use proasic3.all;

entity Cnt4Ref is

    port( Sdram_ctl_v2_0_SD_RefEn : in    std_logic;
          PLL_Test1_0_Sys_66M_Clk : in    std_logic;
          CntEn                   : in    std_logic;
          refenlto5               : out   std_logic
        );

end Cnt4Ref;

architecture DEF_ARCH of Cnt4Ref is 

  component DFN1E1C1
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C1
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AND2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component INV
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component OR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \CntNum[4]\, \CntNum[5]\, \CntNum[3]\, NU_0_1_2, 
        \CntNum[0]\, \CntNum[1]\, XOR2_2_Y, XOR2_3_Y, AND2_2_Y, 
        NU_3_4_5, \CntNum[2]\, INV_0_Y, INV_1_Y, XOR2_0_Y, 
        AND2_1_Y, XOR2_1_Y, AND2_0_Y, \GND\, \VCC\, GND_0, VCC_0
         : std_logic;

begin 


    DFN1E1C1_NU_1 : DFN1E1C1
      port map(D => INV_1_Y, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => Sdram_ctl_v2_0_SD_RefEn, E => CntEn, Q => \CntNum[0]\);
    
    XOR2_1 : XOR2
      port map(A => \CntNum[1]\, B => AND2_0_Y, Y => XOR2_1_Y);
    
    DFN1C1_NU_6 : DFN1C1
      port map(D => XOR2_3_Y, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => Sdram_ctl_v2_0_SD_RefEn, Q => \CntNum[5]\);
    
    AND2_0 : AND2
      port map(A => CntEn, B => \CntNum[0]\, Y => AND2_0_Y);
    
    INV_0 : INV
      port map(A => \CntNum[2]\, Y => INV_0_Y);
    
    DFN1E1C1_NU_5 : DFN1E1C1
      port map(D => XOR2_0_Y, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => Sdram_ctl_v2_0_SD_RefEn, E => NU_0_1_2, Q => 
        \CntNum[4]\);
    
    DFN1C1_NU_2 : DFN1C1
      port map(D => XOR2_1_Y, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => Sdram_ctl_v2_0_SD_RefEn, Q => \CntNum[1]\);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    AND2_1 : AND2
      port map(A => \CntNum[2]\, B => \CntNum[3]\, Y => AND2_1_Y);
    
    XOR2_0 : XOR2
      port map(A => \CntNum[4]\, B => AND2_1_Y, Y => XOR2_0_Y);
    
    XOR2_2 : XOR2
      port map(A => \CntNum[3]\, B => \CntNum[2]\, Y => XOR2_2_Y);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    DFN1C1_NU_6_RNINRGA : OR3C
      port map(A => \CntNum[4]\, B => \CntNum[5]\, C => 
        \CntNum[3]\, Y => refenlto5);
    
    GND_i : GND
      port map(Y => \GND\);
    
    INV_1 : INV
      port map(A => \CntNum[0]\, Y => INV_1_Y);
    
    U_AND3_3_4_5 : AND3
      port map(A => \CntNum[2]\, B => \CntNum[3]\, C => 
        \CntNum[4]\, Y => NU_3_4_5);
    
    XOR2_3 : XOR2
      port map(A => \CntNum[5]\, B => AND2_2_Y, Y => XOR2_3_Y);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    DFN1E1C1_NU_3 : DFN1E1C1
      port map(D => INV_0_Y, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => Sdram_ctl_v2_0_SD_RefEn, E => NU_0_1_2, Q => 
        \CntNum[2]\);
    
    AND2_2 : AND2
      port map(A => NU_0_1_2, B => NU_3_4_5, Y => AND2_2_Y);
    
    DFN1E1C1_NU_4 : DFN1E1C1
      port map(D => XOR2_2_Y, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => Sdram_ctl_v2_0_SD_RefEn, E => NU_0_1_2, Q => 
        \CntNum[3]\);
    
    U_AND3_0_1_2 : AND3
      port map(A => CntEn, B => \CntNum[0]\, C => \CntNum[1]\, Y
         => NU_0_1_2);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3;
use proasic3.all;

entity Counter_ref is

    port( refenlto5               : out   std_logic;
          Sdram_ctl_v2_0_SD_RefEn : in    std_logic;
          PLL_Test1_0_SysRst_O    : in    std_logic;
          PLL_Test1_0_Sys_66M_Clk : in    std_logic;
          Main_ctl4SD_0_ByteRdEn  : in    std_logic;
          CMOS_DrvX_0_LVDSen_2    : in    std_logic
        );

end Counter_ref;

architecture DEF_ARCH of Counter_ref is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component Cnt4Ref
    port( Sdram_ctl_v2_0_SD_RefEn : in    std_logic := 'U';
          PLL_Test1_0_Sys_66M_Clk : in    std_logic := 'U';
          CntEn                   : in    std_logic := 'U';
          refenlto5               : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \CntEn_RNO\, \CntEn\, \GND\, \VCC\, GND_0, VCC_0
         : std_logic;

    for all : Cnt4Ref
	Use entity work.Cnt4Ref(DEF_ARCH);
begin 


    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    CntEn : DFN1C0
      port map(D => \CntEn_RNO\, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \CntEn\);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    CntMap : Cnt4Ref
      port map(Sdram_ctl_v2_0_SD_RefEn => Sdram_ctl_v2_0_SD_RefEn, 
        PLL_Test1_0_Sys_66M_Clk => PLL_Test1_0_Sys_66M_Clk, CntEn
         => \CntEn\, refenlto5 => refenlto5);
    
    CntEn_RNO : NOR2A
      port map(A => CMOS_DrvX_0_LVDSen_2, B => 
        Main_ctl4SD_0_ByteRdEn, Y => \CntEn_RNO\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3;
use proasic3.all;

entity My_adder0_3 is

    port( intData2acc_RNI6J36         : in    std_logic_vector(10 to 10);
          intData2acc_RNIK507         : in    std_logic_vector(9 to 9);
          intData2acc_RNIBJ36         : in    std_logic_vector(15 to 15);
          intData2acc_RNIVOQA         : in    std_logic_vector(0 to 0);
          intData2acc_RNI0TQA         : in    std_logic_vector(1 to 1);
          intData2acc_RNIFHV6         : in    std_logic_vector(4 to 4);
          intData2acc_RNI8J36         : in    std_logic_vector(12 to 12);
          intData2acc_RNIAJ36         : in    std_logic_vector(14 to 14);
          intData2acc_RNI11RA         : in    std_logic_vector(2 to 2);
          intData2acc_RNIEDV6         : in    std_logic_vector(3 to 3);
          intData2acc_RNI9J36         : in    std_logic_vector(13 to 13);
          intData2acc_RNIHPV6         : in    std_logic_vector(6 to 6);
          intData2acc_RNIITV6         : in    std_logic_vector(7 to 7);
          intData2acc_RNI7J36         : in    std_logic_vector(11 to 11);
          intData2acc_RNIDJ36         : in    std_logic_vector(17 to 17);
          intData2acc_RNIGLV6         : in    std_logic_vector(5 to 5);
          intData2acc_RNIJ107         : in    std_logic_vector(8 to 8);
          intData2acc_RNICJ36         : in    std_logic_vector(16 to 16);
          \Z\\My_adder0_0_Sum_[15]\\\ : out   std_logic;
          \Z\\My_adder0_0_Sum_[12]\\\ : out   std_logic;
          \Z\\My_adder0_0_Sum_[6]\\\  : out   std_logic;
          \Z\\My_adder0_0_Sum_[10]\\\ : out   std_logic;
          \Z\\My_adder0_0_Sum_[9]\\\  : out   std_logic;
          \Z\\My_adder0_0_Sum_[7]\\\  : out   std_logic;
          \Z\\My_adder0_0_Sum_[11]\\\ : out   std_logic;
          \Z\\My_adder0_0_Sum_[1]\\\  : out   std_logic;
          \Z\\My_adder0_0_Sum_[3]\\\  : out   std_logic;
          \Z\\My_adder0_0_Sum_[13]\\\ : out   std_logic;
          \Z\\My_adder0_0_Sum_[0]\\\  : out   std_logic;
          \Z\\My_adder0_0_Sum_[8]\\\  : out   std_logic;
          \Z\\My_adder0_0_Sum_[14]\\\ : out   std_logic;
          \Z\\My_adder0_0_Sum_[2]\\\  : out   std_logic;
          \Z\\My_adder0_0_Sum_[4]\\\  : out   std_logic;
          \Z\\My_adder0_0_Sum_[5]\\\  : out   std_logic;
          \Z\\My_adder0_0_Sum_[17]\\\ : out   std_logic;
          My_adder0_3_GND             : in    std_logic;
          \Z\\My_adder0_0_Sum_[16]\\\ : out   std_logic
        );

end My_adder0_3;

architecture DEF_ARCH of My_adder0_3 is 

  component XOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MAJ3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component AND2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal Carry_15_net, Carry_8_net, Carry_7_net, Carry_5_net, 
        Carry_4_net, Carry_16_net, Carry_11_net, Carry_10_net, 
        Carry_6_net, Carry_13_net, Carry_12_net, Carry_3_net, 
        Carry_2_net, Carry_1_net, Carry_14_net, Carry_0_net, 
        Carry_9_net, \GND\, \VCC\, GND_0, VCC_0 : std_logic;

begin 


    XOR3_Sum_16_inst : XOR3
      port map(A => My_adder0_3_GND, B => intData2acc_RNICJ36(16), 
        C => Carry_15_net, Y => \Z\\My_adder0_0_Sum_[16]\\\);
    
    MAJ3_Carry_8_inst : MAJ3
      port map(A => Carry_7_net, B => My_adder0_3_GND, C => 
        intData2acc_RNIJ107(8), Y => Carry_8_net);
    
    MAJ3_Carry_9_inst : MAJ3
      port map(A => Carry_8_net, B => My_adder0_3_GND, C => 
        intData2acc_RNIK507(9), Y => Carry_9_net);
    
    XOR3_Sum_5_inst : XOR3
      port map(A => My_adder0_3_GND, B => intData2acc_RNIGLV6(5), 
        C => Carry_4_net, Y => \Z\\My_adder0_0_Sum_[5]\\\);
    
    XOR3_Sum_2_inst : XOR3
      port map(A => My_adder0_3_GND, B => intData2acc_RNI11RA(2), 
        C => Carry_1_net, Y => \Z\\My_adder0_0_Sum_[2]\\\);
    
    XOR3_Sum_4_inst : XOR3
      port map(A => My_adder0_3_GND, B => intData2acc_RNIFHV6(4), 
        C => Carry_3_net, Y => \Z\\My_adder0_0_Sum_[4]\\\);
    
    XOR3_Sum_11_inst : XOR3
      port map(A => My_adder0_3_GND, B => intData2acc_RNI7J36(11), 
        C => Carry_10_net, Y => \Z\\My_adder0_0_Sum_[11]\\\);
    
    XOR3_Sum_12_inst : XOR3
      port map(A => My_adder0_3_GND, B => intData2acc_RNI8J36(12), 
        C => Carry_11_net, Y => \Z\\My_adder0_0_Sum_[12]\\\);
    
    MAJ3_Carry_5_inst : MAJ3
      port map(A => Carry_4_net, B => My_adder0_3_GND, C => 
        intData2acc_RNIGLV6(5), Y => Carry_5_net);
    
    MAJ3_Carry_2_inst : MAJ3
      port map(A => Carry_1_net, B => My_adder0_3_GND, C => 
        intData2acc_RNI11RA(2), Y => Carry_2_net);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    MAJ3_Carry_1_inst : MAJ3
      port map(A => Carry_0_net, B => My_adder0_3_GND, C => 
        intData2acc_RNI0TQA(1), Y => Carry_1_net);
    
    MAJ3_Carry_4_inst : MAJ3
      port map(A => Carry_3_net, B => My_adder0_3_GND, C => 
        intData2acc_RNIFHV6(4), Y => Carry_4_net);
    
    XOR3_Sum_13_inst : XOR3
      port map(A => My_adder0_3_GND, B => intData2acc_RNI9J36(13), 
        C => Carry_12_net, Y => \Z\\My_adder0_0_Sum_[13]\\\);
    
    XOR3_Sum_1_inst : XOR3
      port map(A => My_adder0_3_GND, B => intData2acc_RNI0TQA(1), 
        C => Carry_0_net, Y => \Z\\My_adder0_0_Sum_[1]\\\);
    
    MAJ3_Carry_12_inst : MAJ3
      port map(A => Carry_11_net, B => My_adder0_3_GND, C => 
        intData2acc_RNI8J36(12), Y => Carry_12_net);
    
    XOR3_Sum_17_inst : XOR3
      port map(A => My_adder0_3_GND, B => intData2acc_RNIDJ36(17), 
        C => Carry_16_net, Y => \Z\\My_adder0_0_Sum_[17]\\\);
    
    MAJ3_Carry_7_inst : MAJ3
      port map(A => Carry_6_net, B => My_adder0_3_GND, C => 
        intData2acc_RNIITV6(7), Y => Carry_7_net);
    
    GND_i : GND
      port map(Y => \GND\);
    
    XOR3_Sum_6_inst : XOR3
      port map(A => My_adder0_3_GND, B => intData2acc_RNIHPV6(6), 
        C => Carry_5_net, Y => \Z\\My_adder0_0_Sum_[6]\\\);
    
    MAJ3_Carry_14_inst : MAJ3
      port map(A => Carry_13_net, B => My_adder0_3_GND, C => 
        intData2acc_RNIAJ36(14), Y => Carry_14_net);
    
    MAJ3_Carry_13_inst : MAJ3
      port map(A => Carry_12_net, B => My_adder0_3_GND, C => 
        intData2acc_RNI9J36(13), Y => Carry_13_net);
    
    XOR3_Sum_3_inst : XOR3
      port map(A => My_adder0_3_GND, B => intData2acc_RNIEDV6(3), 
        C => Carry_2_net, Y => \Z\\My_adder0_0_Sum_[3]\\\);
    
    XOR3_Sum_14_inst : XOR3
      port map(A => My_adder0_3_GND, B => intData2acc_RNIAJ36(14), 
        C => Carry_13_net, Y => \Z\\My_adder0_0_Sum_[14]\\\);
    
    XOR3_Sum_8_inst : XOR3
      port map(A => My_adder0_3_GND, B => intData2acc_RNIJ107(8), 
        C => Carry_7_net, Y => \Z\\My_adder0_0_Sum_[8]\\\);
    
    MAJ3_Carry_11_inst : MAJ3
      port map(A => Carry_10_net, B => My_adder0_3_GND, C => 
        intData2acc_RNI7J36(11), Y => Carry_11_net);
    
    MAJ3_Carry_16_inst : MAJ3
      port map(A => Carry_15_net, B => My_adder0_3_GND, C => 
        intData2acc_RNICJ36(16), Y => Carry_16_net);
    
    XOR3_Sum_7_inst : XOR3
      port map(A => My_adder0_3_GND, B => intData2acc_RNIITV6(7), 
        C => Carry_6_net, Y => \Z\\My_adder0_0_Sum_[7]\\\);
    
    MAJ3_Carry_10_inst : MAJ3
      port map(A => Carry_9_net, B => My_adder0_3_GND, C => 
        intData2acc_RNI6J36(10), Y => Carry_10_net);
    
    MAJ3_Carry_3_inst : MAJ3
      port map(A => Carry_2_net, B => My_adder0_3_GND, C => 
        intData2acc_RNIEDV6(3), Y => Carry_3_net);
    
    XOR3_Sum_15_inst : XOR3
      port map(A => My_adder0_3_GND, B => intData2acc_RNIBJ36(15), 
        C => Carry_14_net, Y => \Z\\My_adder0_0_Sum_[15]\\\);
    
    AND2_Carry_0_inst : AND2
      port map(A => My_adder0_3_GND, B => intData2acc_RNIVOQA(0), 
        Y => Carry_0_net);
    
    MAJ3_Carry_15_inst : MAJ3
      port map(A => Carry_14_net, B => My_adder0_3_GND, C => 
        intData2acc_RNIBJ36(15), Y => Carry_15_net);
    
    XOR3_Sum_9_inst : XOR3
      port map(A => My_adder0_3_GND, B => intData2acc_RNIK507(9), 
        C => Carry_8_net, Y => \Z\\My_adder0_0_Sum_[9]\\\);
    
    XOR2_Sum_0_inst : XOR2
      port map(A => My_adder0_3_GND, B => intData2acc_RNIVOQA(0), 
        Y => \Z\\My_adder0_0_Sum_[0]\\\);
    
    MAJ3_Carry_6_inst : MAJ3
      port map(A => Carry_5_net, B => My_adder0_3_GND, C => 
        intData2acc_RNIHPV6(6), Y => Carry_6_net);
    
    XOR3_Sum_10_inst : XOR3
      port map(A => My_adder0_3_GND, B => intData2acc_RNI6J36(10), 
        C => Carry_9_net, Y => \Z\\My_adder0_0_Sum_[10]\\\);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3;
use proasic3.all;

entity SDRAM_Ref is

    port( \Z\\SDRAM_Ref_0_Ref_state_[2]\\\ : out   std_logic;
          \Z\\SDRAM_Ref_0_Ref_state_[1]\\\ : out   std_logic;
          \Z\\SDRAM_Ref_0_Ref_state_[0]\\\ : out   std_logic;
          ref_ok_1                         : out   std_logic;
          PLL_Test1_0_SysRst_O             : in    std_logic;
          PLL_Test1_0_Sys_66M_Clk          : in    std_logic;
          ref_ok_2                         : out   std_logic;
          Sdram_ctl_v2_0_SD_RefEn          : in    std_logic;
          Sdram_ini_0_Sd_iniOK             : in    std_logic;
          refenlto5                        : in    std_logic;
          Sdram_ctl_v2_0_SD_pdEN           : in    std_logic
        );

end SDRAM_Ref;

architecture DEF_ARCH of SDRAM_Ref is 

  component DFN1E0C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component AO1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AOI1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \DWACT_ADD_CI_0_g_array_1[0]\, 
        \DWACT_ADD_CI_0_TMP[0]\, \SD_refEN_cnt[1]_net_1\, 
        \DWACT_ADD_CI_0_g_array_12[0]\, \SD_refEN_cnt[2]_net_1\, 
        un1_sd_refen_cnt_1, \SD_refEN_cnt[0]_net_1\, 
        un1_sd_refen_cnt_0, \SD_refEN_cnt[3]_net_1\, 
        \pr_state_ns_0[1]\, \pr_state_ns_0_tz[1]\, \un1_refen\, 
        \pr_state[0]_net_1\, \pr_state[5]_net_1\, 
        \pr_state_ns[1]\, \ref_str\, N_101_1, ref_ok_2_0_sqmuxa, 
        \temp[1]_net_1\, ref_ok_1_1_sqmuxa, \pr_state[4]_net_1\, 
        un1_ref_ok_1_1_sqmuxa, \pr_state_RNIVBO[3]_net_1\, 
        \SD_refEN_cnt_4[0]\, \DWACT_ADD_CI_0_partial_sum[0]\, 
        \SD_refEN_cnt_4[3]\, I_17, \temp_4[0]_net_1\, 
        \temp[0]_net_1\, \temp_4[1]_net_1\, \pr_state[3]_net_1\, 
        N_118, \pr_state[2]_net_1\, N_119, \pr_state[1]_net_1\, 
        N_120, \pr_state_RNO_1[2]\, \pr_state_RNO_1[1]\, 
        \pr_state_RNO_0[0]_net_1\, \SD_refEN_cnt_4[1]\, I_15, 
        \SD_refEN_cnt_4[2]\, I_18, \pr_state_RNO[3]_net_1\, N_132, 
        \GND\, \VCC\, GND_0, VCC_0 : std_logic;

begin 


    \Ref_state[0]\ : DFN1E0C0
      port map(D => N_120, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => \pr_state[4]_net_1\, Q => 
        \Z\\SDRAM_Ref_0_Ref_state_[0]\\\);
    
    un1_SD_refEN_cnt_1_I_17 : XOR2
      port map(A => \SD_refEN_cnt[3]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_12[0]\, Y => I_17);
    
    un1_SD_refEN_cnt_1_I_15 : XOR2
      port map(A => \SD_refEN_cnt[1]_net_1\, B => 
        \DWACT_ADD_CI_0_TMP[0]\, Y => I_15);
    
    \pr_state_RNO_0[4]\ : OR2A
      port map(A => \pr_state_ns_0_tz[1]\, B => \un1_refen\, Y
         => \pr_state_ns_0[1]\);
    
    \pr_state_RNO_1[4]\ : AO1
      port map(A => Sdram_ctl_v2_0_SD_pdEN, B => 
        \pr_state[0]_net_1\, C => \pr_state[5]_net_1\, Y => 
        \pr_state_ns_0_tz[1]\);
    
    \temp_4[0]\ : NOR3A
      port map(A => \pr_state[0]_net_1\, B => \temp[1]_net_1\, C
         => \temp[0]_net_1\, Y => \temp_4[0]_net_1\);
    
    \ref_ok_1\ : DFN1C0
      port map(D => ref_ok_1_1_sqmuxa, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => ref_ok_1);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \Ref_state[1]\ : DFN1E0C0
      port map(D => N_119, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => \pr_state[4]_net_1\, Q => 
        \Z\\SDRAM_Ref_0_Ref_state_[1]\\\);
    
    \SD_refEN_cnt_RNI8CH1[3]\ : NOR2A
      port map(A => \SD_refEN_cnt[1]_net_1\, B => 
        \SD_refEN_cnt[3]_net_1\, Y => un1_sd_refen_cnt_0);
    
    \Ref_state[2]\ : DFN1E0C0
      port map(D => \pr_state[0]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => \pr_state[4]_net_1\, Q => 
        \Z\\SDRAM_Ref_0_Ref_state_[2]\\\);
    
    \pr_state[3]\ : DFN1C0
      port map(D => \pr_state_RNO[3]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \pr_state[3]_net_1\);
    
    \SD_refEN_cnt_RNO[0]\ : NOR2B
      port map(A => un1_ref_ok_1_1_sqmuxa, B => 
        \DWACT_ADD_CI_0_partial_sum[0]\, Y => \SD_refEN_cnt_4[0]\);
    
    \SD_refEN_cnt_RNO[1]\ : MX2
      port map(A => \pr_state[4]_net_1\, B => I_15, S => 
        un1_ref_ok_1_1_sqmuxa, Y => \SD_refEN_cnt_4[1]\);
    
    \pr_state_RNO_0[0]\ : AO1A
      port map(A => Sdram_ctl_v2_0_SD_pdEN, B => 
        \pr_state[0]_net_1\, C => \pr_state[2]_net_1\, Y => N_118);
    
    \SD_refEN_cnt[3]\ : DFN1C0
      port map(D => \SD_refEN_cnt_4[3]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \SD_refEN_cnt[3]_net_1\);
    
    \temp[1]\ : DFN1C0
      port map(D => \temp_4[1]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \temp[1]_net_1\);
    
    \SD_refEN_cnt_RNI6CH1[0]\ : NOR2A
      port map(A => \SD_refEN_cnt[2]_net_1\, B => 
        \SD_refEN_cnt[0]_net_1\, Y => un1_sd_refen_cnt_1);
    
    \pr_state[2]\ : DFN1C0
      port map(D => \pr_state_RNO_1[2]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \pr_state[2]_net_1\);
    
    un1_SD_refEN_cnt_1_I_19 : NOR2B
      port map(A => \DWACT_ADD_CI_0_TMP[0]\, B => 
        \SD_refEN_cnt[1]_net_1\, Y => 
        \DWACT_ADD_CI_0_g_array_1[0]\);
    
    \pr_state_RNO[0]\ : NOR2A
      port map(A => N_118, B => \un1_refen\, Y => 
        \pr_state_RNO_0[0]_net_1\);
    
    ref_str : DFN1E0C0
      port map(D => \pr_state[4]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => un1_ref_ok_1_1_sqmuxa, Q => \ref_str\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \SD_refEN_cnt[1]\ : DFN1C0
      port map(D => \SD_refEN_cnt_4[1]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \SD_refEN_cnt[1]_net_1\);
    
    \pr_state_RNO[4]\ : AO1C
      port map(A => \ref_str\, B => N_101_1, C => 
        \pr_state_ns_0[1]\, Y => \pr_state_ns[1]\);
    
    \pr_state_RNO[1]\ : NOR2A
      port map(A => \pr_state[3]_net_1\, B => \un1_refen\, Y => 
        \pr_state_RNO_1[1]\);
    
    \pr_state[0]\ : DFN1C0
      port map(D => \pr_state_RNO_0[0]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \pr_state[0]_net_1\);
    
    \pr_state_RNO[2]\ : NOR2A
      port map(A => \pr_state[1]_net_1\, B => \un1_refen\, Y => 
        \pr_state_RNO_1[2]\);
    
    un1_SD_refEN_cnt_1_I_21 : NOR2B
      port map(A => \DWACT_ADD_CI_0_g_array_1[0]\, B => 
        \SD_refEN_cnt[2]_net_1\, Y => 
        \DWACT_ADD_CI_0_g_array_12[0]\);
    
    un1_SD_refEN_cnt_1_I_11 : XOR2
      port map(A => \SD_refEN_cnt[0]_net_1\, B => 
        \pr_state_RNIVBO[3]_net_1\, Y => 
        \DWACT_ADD_CI_0_partial_sum[0]\);
    
    \temp[0]\ : DFN1C0
      port map(D => \temp_4[0]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \temp[0]_net_1\);
    
    \pr_state_RNIVBO[3]\ : OR2
      port map(A => \pr_state[4]_net_1\, B => \pr_state[3]_net_1\, 
        Y => \pr_state_RNIVBO[3]_net_1\);
    
    un1_SD_refEN_cnt_1_I_1 : AND2
      port map(A => \SD_refEN_cnt[0]_net_1\, B => 
        \pr_state_RNIVBO[3]_net_1\, Y => \DWACT_ADD_CI_0_TMP[0]\);
    
    \pr_state[4]\ : DFN1C0
      port map(D => \pr_state_ns[1]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \pr_state[4]_net_1\);
    
    un2_sd_refen : OR2B
      port map(A => Sdram_ini_0_Sd_iniOK, B => 
        Sdram_ctl_v2_0_SD_RefEn, Y => N_132);
    
    ref_ok_2_RNO : NOR2B
      port map(A => \temp[1]_net_1\, B => \pr_state[0]_net_1\, Y
         => ref_ok_2_0_sqmuxa);
    
    \pr_state_RNIJ9OK[4]\ : NOR2A
      port map(A => \pr_state[4]_net_1\, B => \un1_refen\, Y => 
        N_101_1);
    
    \temp_4[1]\ : NOR3B
      port map(A => \pr_state[0]_net_1\, B => \temp[0]_net_1\, C
         => \temp[1]_net_1\, Y => \temp_4[1]_net_1\);
    
    \Ref_state_RNO[0]\ : OR2
      port map(A => \pr_state[3]_net_1\, B => \pr_state[2]_net_1\, 
        Y => N_120);
    
    \ref_ok_2\ : DFN1C0
      port map(D => ref_ok_2_0_sqmuxa, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => ref_ok_2);
    
    \pr_state[1]\ : DFN1C0
      port map(D => \pr_state_RNO_1[1]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \pr_state[1]_net_1\);
    
    \SD_refEN_cnt[0]\ : DFN1C0
      port map(D => \SD_refEN_cnt_4[0]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \SD_refEN_cnt[0]_net_1\);
    
    \pr_state[5]\ : DFN1P0
      port map(D => \un1_refen\, CLK => PLL_Test1_0_Sys_66M_Clk, 
        PRE => PLL_Test1_0_SysRst_O, Q => \pr_state[5]_net_1\);
    
    un1_refen : NOR2B
      port map(A => N_132, B => refenlto5, Y => \un1_refen\);
    
    \SD_refEN_cnt_RNO[2]\ : MX2
      port map(A => \pr_state[4]_net_1\, B => I_18, S => 
        un1_ref_ok_1_1_sqmuxa, Y => \SD_refEN_cnt_4[2]\);
    
    \pr_state_RNIEUE3[4]\ : AOI1B
      port map(A => un1_sd_refen_cnt_1, B => un1_sd_refen_cnt_0, 
        C => \pr_state[4]_net_1\, Y => ref_ok_1_1_sqmuxa);
    
    un1_SD_refEN_cnt_1_I_18 : XOR2
      port map(A => \SD_refEN_cnt[2]_net_1\, B => 
        \DWACT_ADD_CI_0_g_array_1[0]\, Y => I_18);
    
    \pr_state_RNIDA74[4]\ : OR2A
      port map(A => \pr_state_RNIVBO[3]_net_1\, B => 
        ref_ok_1_1_sqmuxa, Y => un1_ref_ok_1_1_sqmuxa);
    
    \SD_refEN_cnt_RNO[3]\ : NOR2B
      port map(A => un1_ref_ok_1_1_sqmuxa, B => I_17, Y => 
        \SD_refEN_cnt_4[3]\);
    
    \pr_state_RNO[3]\ : NOR2B
      port map(A => \ref_str\, B => N_101_1, Y => 
        \pr_state_RNO[3]_net_1\);
    
    \SD_refEN_cnt[2]\ : DFN1C0
      port map(D => \SD_refEN_cnt_4[2]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \SD_refEN_cnt[2]_net_1\);
    
    \Ref_state_RNO[1]\ : OR2
      port map(A => \pr_state[2]_net_1\, B => \pr_state[1]_net_1\, 
        Y => N_119);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3;
use proasic3.all;

entity WaveGenSingleZ18 is

    port( Sdram_cmd_0_RFifo_we    : out   std_logic;
          PLL_Test1_0_SysRst_O    : in    std_logic;
          PLL_Test1_0_Sys_66M_Clk : in    std_logic;
          Rfifo_weEN              : in    std_logic
        );

end WaveGenSingleZ18;

architecture DEF_ARCH of WaveGenSingleZ18 is 

  component INV
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component OR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal Rfifo_weEN_i, N_106, \PrState[1]_net_1\, 
        \Phase2Cnt[0]_net_1\, \Phase1Cnt_RNO_3[2]\, N_93, 
        \Phase1Cnt[2]_net_1\, \PrState[2]_net_1\, 
        \Phase1Cnt_RNO_1[1]\, \Phase1Cnt[0]_net_1\, 
        \Phase1Cnt[1]_net_1\, \PrState_ns_0_tz[2]\, N_94, 
        \CycCnt[0]_net_1\, \DelayCnt_RNIS6G6[0]_net_1\, 
        \PrState_ns[2]\, N_103, N_107_1, N_95, 
        \PrState_RNO_0_0[3]\, \PrState[3]_net_1\, 
        \DelayCnt[0]_net_1\, \CycCnt_RNO_5[0]\, 
        \PrState[4]_net_1\, \PrState_ns[3]\, N_85_i_0, 
        Phase1Cnt_n0, \GND\, \VCC\, GND_0, VCC_0 : std_logic;

begin 


    \PrState_RNO[4]\ : INV
      port map(A => Rfifo_weEN, Y => Rfifo_weEN_i);
    
    \PrState_RNO[2]\ : AO1B
      port map(A => \PrState_ns_0_tz[2]\, B => Rfifo_weEN, C => 
        N_103, Y => \PrState_ns[2]\);
    
    \DelayCnt[0]\ : DFN1C0
      port map(D => \DelayCnt_RNIS6G6[0]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \DelayCnt[0]_net_1\);
    
    \PrState_RNI5AU7[2]\ : NOR2B
      port map(A => \PrState[2]_net_1\, B => Rfifo_weEN, Y => 
        N_107_1);
    
    WFO : DFN1C0
      port map(D => \PrState[2]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => Sdram_cmd_0_RFifo_we);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    \PrState[3]\ : DFN1C0
      port map(D => N_85_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \PrState[3]_net_1\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \PrState[1]\ : DFN1C0
      port map(D => \PrState_ns[3]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \PrState[1]_net_1\);
    
    \PrState_RNO_0[1]\ : OR3C
      port map(A => \PrState[1]_net_1\, B => \Phase2Cnt[0]_net_1\, 
        C => Rfifo_weEN, Y => N_106);
    
    \CycCnt[0]\ : DFN1C0
      port map(D => \CycCnt_RNO_5[0]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \CycCnt[0]_net_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \PrState_RNO[1]\ : AO1C
      port map(A => N_95, B => N_107_1, C => N_106, Y => 
        \PrState_ns[3]\);
    
    \Phase1Cnt[1]\ : DFN1C0
      port map(D => \Phase1Cnt_RNO_1[1]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \Phase1Cnt[1]_net_1\);
    
    \PrState_RNO[3]\ : OA1
      port map(A => \PrState_RNO_0_0[3]\, B => \PrState[4]_net_1\, 
        C => Rfifo_weEN, Y => N_85_i_0);
    
    \PrState[4]\ : DFN1P0
      port map(D => Rfifo_weEN_i, CLK => PLL_Test1_0_Sys_66M_Clk, 
        PRE => PLL_Test1_0_SysRst_O, Q => \PrState[4]_net_1\);
    
    \Phase1Cnt_RNO[0]\ : NOR2A
      port map(A => \PrState[2]_net_1\, B => \Phase1Cnt[0]_net_1\, 
        Y => Phase1Cnt_n0);
    
    \Phase1Cnt_RNIBBBE[2]\ : OR2B
      port map(A => \Phase1Cnt[2]_net_1\, B => N_93, Y => N_95);
    
    \CycCnt_RNO[0]\ : XA1B
      port map(A => \CycCnt[0]_net_1\, B => N_94, C => 
        \PrState[4]_net_1\, Y => \CycCnt_RNO_5[0]\);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    \Phase1Cnt_RNO[1]\ : XA1
      port map(A => \Phase1Cnt[0]_net_1\, B => 
        \Phase1Cnt[1]_net_1\, C => \PrState[2]_net_1\, Y => 
        \Phase1Cnt_RNO_1[1]\);
    
    \Phase1Cnt_RNO[2]\ : XA1
      port map(A => N_93, B => \Phase1Cnt[2]_net_1\, C => 
        \PrState[2]_net_1\, Y => \Phase1Cnt_RNO_3[2]\);
    
    \Phase1Cnt_RNIH7I9[1]\ : NOR2B
      port map(A => \Phase1Cnt[1]_net_1\, B => 
        \Phase1Cnt[0]_net_1\, Y => N_93);
    
    \PrState_RNO_1[2]\ : OR2B
      port map(A => N_107_1, B => N_95, Y => N_103);
    
    \Phase1Cnt[0]\ : DFN1C0
      port map(D => Phase1Cnt_n0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[0]_net_1\);
    
    \Phase2Cnt_RNI2Q7A[0]\ : NOR2A
      port map(A => \PrState[1]_net_1\, B => \Phase2Cnt[0]_net_1\, 
        Y => N_94);
    
    \Phase2Cnt[0]\ : DFN1C0
      port map(D => N_94, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase2Cnt[0]_net_1\);
    
    \PrState_RNO_0[2]\ : AO1
      port map(A => N_94, B => \CycCnt[0]_net_1\, C => 
        \DelayCnt_RNIS6G6[0]_net_1\, Y => \PrState_ns_0_tz[2]\);
    
    \Phase1Cnt[2]\ : DFN1C0
      port map(D => \Phase1Cnt_RNO_3[2]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \Phase1Cnt[2]_net_1\);
    
    \PrState_RNO_0[3]\ : NOR2B
      port map(A => \PrState[3]_net_1\, B => \DelayCnt[0]_net_1\, 
        Y => \PrState_RNO_0_0[3]\);
    
    \PrState[2]\ : DFN1C0
      port map(D => \PrState_ns[2]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \PrState[2]_net_1\);
    
    \DelayCnt_RNIS6G6[0]\ : NOR2A
      port map(A => \PrState[3]_net_1\, B => \DelayCnt[0]_net_1\, 
        Y => \DelayCnt_RNIS6G6[0]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3;
use proasic3.all;

entity Sdram_cmd is

    port( SD_cs_n_c_c                      : out   std_logic_vector(1 to 1);
          SD_dqm_c_c_c_c_c_c_c_c           : out   std_logic_vector(1 to 1);
          SD_cke_c_c                       : in    std_logic_vector(0 to 0);
          SD_Clk_c_c                       : out   std_logic_vector(1 to 1);
          SD_addr_c                        : out   std_logic_vector(12 downto 0);
          Sdram_cmd_0_RFifo_we             : out   std_logic;
          Sdram_cmd_0_rdrow_end            : out   std_logic;
          Sdram_cmd_0_WFifo_re             : out   std_logic;
          Sdram_cmd_0_wrrow_end            : out   std_logic;
          SD_ras_n_c                       : out   std_logic;
          SD_we_n_c                        : out   std_logic;
          SD_cas_n_c                       : out   std_logic;
          CMOS_DrvX_0_LVDSen               : in    std_logic;
          Sdram_cmd_0_SDoneFrameOk         : out   std_logic;
          CMOS_DrvX_0_SDramEn              : in    std_logic;
          PLL_Test1_0_SysRst_O             : in    std_logic;
          PLL_Test1_0_Sys_66M_Clk          : in    std_logic;
          LVDS_enReg                       : out   std_logic;
          CMOS_DrvX_0_LVDSen_2             : in    std_logic;
          \Z\\Sdram_ini_0_ini_state_[0]\\\ : in    std_logic;
          un6_sdramenreg                   : in    std_logic;
          N_264                            : out   std_logic;
          \Z\\SDRAM_Ref_0_Ref_state_[0]\\\ : in    std_logic;
          \Z\\SDRAM_Ref_0_Ref_state_[2]\\\ : in    std_logic;
          \Z\\SDRAM_Ref_0_Ref_state_[1]\\\ : in    std_logic;
          PLL_Test1_0_Sdram_clk            : in    std_logic;
          \Z\\SDram_rd_0_rd_state_[1]\\\   : in    std_logic;
          \Z\\SDram_rd_0_rd_state_[2]\\\   : in    std_logic;
          \Z\\SDram_rd_0_rd_state_[0]\\\   : in    std_logic;
          \Z\\Sdram_ini_0_ini_state_[2]\\\ : in    std_logic;
          \Z\\Sdram_ini_0_ini_state_[1]\\\ : in    std_logic;
          N_264_0                          : out   std_logic;
          N_264_1                          : out   std_logic;
          \Z\\SDRAM_wr_0_wr_state_[1]\\\   : in    std_logic;
          \Z\\SDRAM_wr_0_wr_state_[0]\\\   : in    std_logic;
          \Z\\SDRAM_wr_0_wr_state_[2]\\\   : in    std_logic;
          N_264_2                          : out   std_logic
        );

end Sdram_cmd;

architecture DEF_ARCH of Sdram_cmd is 

  component OR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NOR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component XA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OAI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XO1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1E
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E0C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MX2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E1
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component XNOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component WaveGenSingleZ18
    port( Sdram_cmd_0_RFifo_we    : out   std_logic;
          PLL_Test1_0_SysRst_O    : in    std_logic := 'U';
          PLL_Test1_0_Sys_66M_Clk : in    std_logic := 'U';
          Rfifo_weEN              : in    std_logic := 'U'
        );
  end component;

  component MX2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal N_186_0, ADD_13x13_medium_area_I48_Y_0_0, 
        \SD_wrAddr_row[11]_net_1\, sd_wraddr_row20, 
        ADD_13x13_medium_area_I49_Y_0_0, 
        \SD_wrAddr_row[12]_net_1\, 
        ADD_13x13_medium_area_I47_Y_0_0, 
        \SD_wrAddr_row[10]_net_1\, 
        ADD_13x13_medium_area_I22_un1_Y_1, N242, 
        ADD_13x13_medium_area_I15_Y_1, \SD_wrAddr_row[6]_net_1\, 
        \SD_wrAddr_row[7]_net_1\, N253, 
        ADD_13x13_medium_area_I48_Y_0_0_0, 
        \SD_rdAddr_row[11]_net_1\, sd_rdaddr_row18_i, 
        \addr_11_0_i_2[6]\, \addr_RNO_2[6]_net_1\, 
        \addr_RNO_3[6]_net_1\, \addr_RNO_4[6]_net_1\, 
        \addr_11_0_i_1[6]\, N_191, \addr_RNO_5[6]_net_1\, 
        \addr_11_0_i_2[4]\, \addr_RNO_2[4]_net_1\, 
        \addr_RNO_3[4]_net_1\, \addr_RNO_4[4]_net_1\, 
        \addr_11_0_i_1[4]\, \SD_wrAddr_row[4]_net_1\, 
        \addr_RNO_5[4]_net_1\, \addr_11_0_i_2[3]\, 
        \addr_RNO_2[3]_net_1\, \addr_RNO_3[3]_net_1\, 
        \addr_11_0_i_0[3]\, N_372, \SD_WrAddr_col[3]_net_1\, 
        \addr_RNO_5[3]_net_1\, \addr_11_i_i_2[5]\, N_319, N_323, 
        N_322, \addr_11_i_i_1[5]\, \SD_wrAddr_row[5]_net_1\, 
        N_320, \addr_11_0_i_2[7]\, \addr_RNO_2[7]_net_1\, N_333, 
        \addr_RNO_4[7]_net_1\, \addr_11_0_i_1[7]\, N_331, 
        \addr_11_0_i_2[8]\, \addr_RNO_2[8]_net_1\, N_338, 
        \addr_RNO_4[8]_net_1\, \addr_11_0_i_1[8]\, 
        \SD_wrAddr_row[8]_net_1\, N_336, \addr_11_i_0_2[9]\, 
        \addr_RNO_2[9]_net_1\, N_253, \addr_RNO_4[9]_net_1\, 
        \addr_11_i_0_1[9]\, \SD_wrAddr_row[9]_net_1\, N_251, 
        \addr_11_0_0_0[1]\, \SD_wrAddr_row[1]_net_1\, N_303, 
        \addr_11_0_0_0[0]\, \SD_wrAddr_row[0]_net_1\, N_300, 
        ADD_13x13_medium_area_I49_Y_0_0_0, 
        \SD_rdAddr_row[12]_net_1\, ADD_13x13_medium_area_I14_Y_0, 
        \SD_wrAddr_row[3]_net_1\, \SD_wrAddr_row[2]_net_1\, 
        we_n_4_0_0_1, \we_n_RNO_2\, N_362, N_360, 
        \addr_11_0_i_2[2]\, N_371, \addr_RNO_4[2]_net_1\, 
        \addr_11_0_i_0[2]\, \addr_11_0_i_a7_0[2]\, N_192, N_308, 
        ras_n_5_7_0_0_0, N_221, N_187, N_635, 
        ADD_13x13_medium_area_I22_un1_Y_1_0, 
        ADD_13x13_medium_area_I22_un1_Y_0, N199, N242_0, 
        \addr_14_i_0_3[10]\, N_365, N_366, \addr_14_i_0_1[10]\, 
        N_367, \addr_RNO_7[10]_net_1\, N_364, cas_n_4_6_0_0_1, 
        N_637, N_241, N_638, \cs_n_5_0_iv_0_0_1[0]\, N_358, 
        \cs_n_1_RNO_4[0]_net_1\, N_355, 
        ADD_13x13_medium_area_I15_Y_1_0, \SD_rdAddr_row[6]_net_1\, 
        \SD_rdAddr_row[7]_net_1\, N253_0, cas_n_4_6_0_a7_1_0, 
        N_384, \un1_sd_wraddr_row8_i_1[12]\, 
        \un1_sd_wraddr_row8_i_0[12]\, N_239, 
        \SD_WrAddr_col[10]_net_1\, N_238, 
        ADD_13x13_medium_area_I14_Y_0_0, \SD_rdAddr_row[3]_net_1\, 
        \SD_rdAddr_row[2]_net_1\, un1_cs_n7_4_i_0_a7_1, 
        un1_cs_n7_4_i_0_a7_0, \temp_w[3]_net_1\, 
        sd_wraddr_row20_0_a7_9, sd_wraddr_row20_0_a7_6, 
        sd_wraddr_row20_0_a7_8, sd_wraddr_row20_0_a7_4, 
        sd_wraddr_row20_0_a7_7, sd_wraddr_row20_0_a7_2, 
        sd_rdaddr_row18_0_a7_9, sd_rdaddr_row18_0_a7_6, 
        \SD_rdAddr_row[4]_net_1\, sd_rdaddr_row18_0_a7_8, 
        sd_rdaddr_row18_0_a7_4, \SD_rdAddr_row[5]_net_1\, 
        sd_rdaddr_row18_0_a7_7, sd_rdaddr_row18_0_a7_2, 
        \SD_rdAddr_row[1]_net_1\, \SD_rdAddr_row[0]_net_1\, 
        \SD_rdAddr_row[10]_net_1\, \SD_rdAddr_row[8]_net_1\, 
        \SD_rdAddr_row[9]_net_1\, un4lt10_i_a2_0_a7_3, 
        \SD_rdAddr_col[5]_net_1\, \SD_rdAddr_col[4]_net_1\, 
        \SD_rdAddr_col[10]_net_1\, un4lt10_i_a2_0_a7_2, 
        \SD_rdAddr_col[8]_net_1\, \SD_rdAddr_col[9]_net_1\, 
        un4lt10_i_a2_0_a7_1, \SD_rdAddr_col[6]_net_1\, 
        \SD_rdAddr_col[7]_net_1\, \un1_sd_wraddr_row8_i_o7_1[12]\, 
        \SD_WrAddr_col[7]_net_1\, \SD_WrAddr_col[8]_net_1\, 
        \un1_sd_wraddr_row8_i_o7_0[12]\, \SD_WrAddr_col[5]_net_1\, 
        \SD_WrAddr_col[6]_net_1\, \temp_w_n1_0_i_0\, 
        \temp_w[0]_net_1\, \temp_w[1]_net_1\, \temp_w_n2_0_i_0\, 
        N_207, \temp_w[2]_net_1\, N_12_i_0, we_n_4, N_216, N_361, 
        \cs_n_5[0]\, N_357, N_356, N_6_i_0, N_249_i, N_190, N_211, 
        N_223, N_224, N_193, N_198, N_370, N_205, N_174_i_0, 
        N_248, N_261, SD_WrAddr_cole, un7_sdram_enreg, N_7, N_19, 
        N_209, \SD_WrAddr_col[9]_net_1\, un1_sdram_enreg_2, N_17, 
        N_203, N_15, N_199, N_13, N_196, ras_n_5, N_634, N_542, 
        N_204, N_297, N_428, N_543, N_544, N_214, N_565, N_541, 
        N_197, N_35, N_195, N_540, \SD_rdAddr_col[3]_net_1\, 
        N_178, N_343, N_345, N_344, N_172_i_0, N245, N256, N215, 
        N_189, N_383, \dqm_1_RNO[0]_net_1\, N_263, \N_264_0\, 
        N_168, cas_n_4, N_353_2, N_220, \addr_11[0]\, N_630, 
        \addr_11[1]\, N_304, N_9_i_0, \SD_WrAddr_col[4]_net_1\, 
        N_11_i_0, N_255, N_164_i_0, \addr_RNO_1[3]_net_1\, N_633, 
        N_176, N_340, N_342, N_162_i_0, N_166_i_0, N_170_i_0, 
        N245_0, N256_0, N215_0, N153, I34_un1_Y, 
        \SD_wrAddr_row_6[0]\, \SD_wrAddr_row_6[9]\, N_225, N_10, 
        N_217, \temp_w_n0_0_i_0\, \temp_w_n3_0_i_0\, 
        \SD_wrAddr_row_6[8]\, N_21, N_218, N_4, N_186, N_201, 
        N_202, N_219, SD_rdAddr_cole, SD_rdAddr_col_n0, 
        \SD_rdAddr_col_RNO[10]_net_1\, N261, N247, 
        \un1_SD_rdAddr_row_i[1]\, \SD_rdAddr_row_6[0]\, N_539, 
        \SD_rdAddr_row_6[1]\, \SD_rdAddr_row_6[10]\, 
        \SD_rdAddr_row_6[11]\, N_343_1, \SD_rdAddr_row_6[12]\, 
        N237, \SD_rdAddr_row_6[9]\, I34_un1_Y_0, 
        \SD_rdAddr_row_6[8]\, \SD_rdAddr_row_6[7]\, I35_un1_Y, 
        \SD_rdAddr_row_6[6]\, N258, \SD_rdAddr_row_6[5]\, 
        I36_un1_Y, \SD_rdAddr_row_6[4]\, \SD_rdAddr_row_6[3]\, 
        I37_un1_Y, \SD_rdAddr_row_6[2]\, un1_rfifo_ween2_3, 
        \Rfifo_weEN\, N_231, N237_0, N247_0, N261_i, 
        \SD_wrAddr_row_6[10]\, \SD_wrAddr_row_6[11]\, 
        \SD_wrAddr_row_6[12]\, N_379, \SD_wrAddr_row_6[5]\, 
        I36_un1_Y_0, N_16, \SD_wrAddr_row_6[7]\, I35_un1_Y_0, 
        \SD_wrAddr_row_6[6]\, N258_0, \SD_wrAddr_row_6[4]\, 
        \SD_wrAddr_row_6[3]\, I37_un1_Y_0, \SD_wrAddr_row_6[2]\, 
        \SD_wrAddr_row_6[1]\, \sdram_enReg\, \dly3_SDoneFrameOk\, 
        \dly2_SDoneFrameOk\, \dly1_SDoneFrameOk\, \SD_addr_c[0]\, 
        \SD_addr_c[1]\, \SD_addr_c[2]\, \SD_addr_c[3]\, 
        \SD_addr_c[4]\, \SD_addr_c[5]\, \SD_addr_c[6]\, 
        \SD_addr_c[7]\, \SD_addr_c[8]\, \SD_addr_c[9]\, 
        \SD_addr_c[10]\, \SD_addr_c[11]\, \SD_addr_c[12]\, \GND\, 
        \VCC\, GND_0, VCC_0 : std_logic;

    for all : WaveGenSingleZ18
	Use entity work.WaveGenSingleZ18(DEF_ARCH);
begin 

    SD_addr_c(12) <= \SD_addr_c[12]\;
    SD_addr_c(11) <= \SD_addr_c[11]\;
    SD_addr_c(10) <= \SD_addr_c[10]\;
    SD_addr_c(9) <= \SD_addr_c[9]\;
    SD_addr_c(8) <= \SD_addr_c[8]\;
    SD_addr_c(7) <= \SD_addr_c[7]\;
    SD_addr_c(6) <= \SD_addr_c[6]\;
    SD_addr_c(5) <= \SD_addr_c[5]\;
    SD_addr_c(4) <= \SD_addr_c[4]\;
    SD_addr_c(3) <= \SD_addr_c[3]\;
    SD_addr_c(2) <= \SD_addr_c[2]\;
    SD_addr_c(1) <= \SD_addr_c[1]\;
    SD_addr_c(0) <= \SD_addr_c[0]\;
    N_264_0 <= \N_264_0\;

    \addr_RNO_2[4]\ : OR3A
      port map(A => N_186, B => N_189, C => \SD_addr_c[4]\, Y => 
        \addr_RNO_2[4]_net_1\);
    
    un1_rfifo_ween2_3_0_0_o4_0 : NOR2A
      port map(A => \Z\\SDram_rd_0_rd_state_[0]\\\, B => 
        \Z\\SDram_rd_0_rd_state_[2]\\\, Y => N_220);
    
    \cs_n_1_RNO_0[0]\ : NOR3C
      port map(A => N_358, B => \cs_n_1_RNO_4[0]_net_1\, C => 
        N_355, Y => \cs_n_5_0_iv_0_0_1[0]\);
    
    \addr_RNO_1[7]\ : OA1
      port map(A => N_191, B => \SD_wrAddr_row[7]_net_1\, C => 
        N_331, Y => \addr_11_0_i_1[7]\);
    
    ras_n_RNO : OR3C
      port map(A => N_634, B => ras_n_5_7_0_0_0, C => N_216, Y
         => ras_n_5);
    
    \addr[11]\ : DFN1C0
      port map(D => N_176, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \SD_addr_c[11]\);
    
    we_n_RNO_3 : OR2A
      port map(A => \Z\\SDRAM_Ref_0_Ref_state_[1]\\\, B => N_187, 
        Y => N_362);
    
    \addr_RNO_3[8]\ : OR2
      port map(A => \SD_WrAddr_col[8]_net_1\, B => N_372, Y => 
        N_338);
    
    \SD_rdAddr_row[2]\ : DFN1C0
      port map(D => \SD_rdAddr_row_6[2]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \SD_rdAddr_row[2]_net_1\);
    
    \addr_11_i_0_a7[9]\ : OR3A
      port map(A => N_186, B => N_189, C => N_384, Y => N_249_i);
    
    \SD_rdAddr_row[3]\ : DFN1C0
      port map(D => \SD_rdAddr_row_6[3]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \SD_rdAddr_row[3]_net_1\);
    
    \cs_n_1[0]\ : DFN1P0
      port map(D => \cs_n_5[0]\, CLK => PLL_Test1_0_Sys_66M_Clk, 
        PRE => PLL_Test1_0_SysRst_O, Q => SD_cs_n_c_c(1));
    
    cas_n_RNO_1 : NOR3C
      port map(A => N_637, B => N_241, C => N_638, Y => 
        cas_n_4_6_0_0_1);
    
    \addr[7]\ : DFN1C0
      port map(D => N_172_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \SD_addr_c[7]\);
    
    \SD_rdAddr_row_RNIQAP2[1]\ : NOR3A
      port map(A => sd_rdaddr_row18_0_a7_2, B => 
        \SD_rdAddr_row[1]_net_1\, C => \SD_rdAddr_row[0]_net_1\, 
        Y => sd_rdaddr_row18_0_a7_7);
    
    \SD_WrAddr_col_RNI9IMM[8]\ : NOR2B
      port map(A => \SD_WrAddr_col[8]_net_1\, B => N_203, Y => 
        N_209);
    
    \SD_rdAddr_col[6]\ : DFN1E1C0
      port map(D => N_541, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => SD_rdAddr_cole, Q => 
        \SD_rdAddr_col[6]_net_1\);
    
    \SD_wrAddr_row_RNO[7]\ : XA1A
      port map(A => \SD_wrAddr_row[7]_net_1\, B => I35_un1_Y_0, C
         => un7_sdram_enreg, Y => \SD_wrAddr_row_6[7]\);
    
    \SD_wrAddr_row_RNIRNGQ[4]\ : NOR3A
      port map(A => sd_wraddr_row20_0_a7_6, B => 
        \SD_wrAddr_row[6]_net_1\, C => \SD_wrAddr_row[4]_net_1\, 
        Y => sd_wraddr_row20_0_a7_9);
    
    Rfifo_weEN_RNO : AO1
      port map(A => \Rfifo_weEN\, B => N_205, C => N_220, Y => 
        un1_rfifo_ween2_3);
    
    \dqm_4_iv_i_0_a7_0_0[0]\ : NOR3A
      port map(A => \Z\\SDRAM_wr_0_wr_state_[2]\\\, B => 
        \Z\\SDRAM_wr_0_wr_state_[0]\\\, C => 
        \Z\\SDRAM_wr_0_wr_state_[1]\\\, Y => \N_264_0\);
    
    \addr_RNO_4[8]\ : OR3A
      port map(A => N_186_0, B => N_371, C => 
        \SD_rdAddr_col[8]_net_1\, Y => \addr_RNO_4[8]_net_1\);
    
    \SD_rdAddr_row[12]\ : DFN1C0
      port map(D => \SD_rdAddr_row_6[12]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \SD_rdAddr_row[12]_net_1\);
    
    \SD_rdAddr_col[3]\ : DFN1E1C0
      port map(D => SD_rdAddr_col_n0, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => SD_rdAddr_cole, Q => \SD_rdAddr_col[3]_net_1\);
    
    \dqm_1_RNO[0]\ : NOR3A
      port map(A => N_372, B => N_263, C => \N_264_0\, Y => 
        \dqm_1_RNO[0]_net_1\);
    
    \addr_RNO_2[11]\ : NOR3A
      port map(A => N_191, B => N_192, C => 
        \SD_rdAddr_row[11]_net_1\, Y => N_633);
    
    \addr_RNO_4[2]\ : OR3A
      port map(A => N_186, B => N_192, C => 
        \SD_rdAddr_row[2]_net_1\, Y => \addr_RNO_4[2]_net_1\);
    
    \addr_RNO[5]\ : OR3C
      port map(A => \addr_11_i_i_2[5]\, B => \addr_11_i_i_1[5]\, 
        C => N_249_i, Y => N_168);
    
    \SD_wrAddr_row_RNO[8]\ : XA1
      port map(A => \SD_wrAddr_row[8]_net_1\, B => N245_0, C => 
        un7_sdram_enreg, Y => \SD_wrAddr_row_6[8]\);
    
    \SD_WrAddr_col_RNO[6]\ : XA1C
      port map(A => N_196, B => \SD_WrAddr_col[6]_net_1\, C => 
        un1_sdram_enreg_2, Y => N_13);
    
    \SD_rdAddr_row[7]\ : DFN1C0
      port map(D => \SD_rdAddr_row_6[7]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \SD_rdAddr_row[7]_net_1\);
    
    sdram_enReg_RNIU39L : OR2A
      port map(A => un7_sdram_enreg, B => un6_sdramenreg, Y => 
        N_202);
    
    \addr_RNO_3[7]\ : OR2
      port map(A => \SD_WrAddr_col[7]_net_1\, B => N_372, Y => 
        N_333);
    
    \addr_RNO_0[0]\ : OA1A
      port map(A => \SD_wrAddr_row[0]_net_1\, B => N_191, C => 
        N_300, Y => \addr_11_0_0_0[0]\);
    
    \addr_RNO_2[9]\ : OR3A
      port map(A => N_186_0, B => N_189, C => \SD_addr_c[9]\, Y
         => \addr_RNO_2[9]_net_1\);
    
    ras_n_5_7_0_a2_3 : OR2B
      port map(A => \Z\\SDram_rd_0_rd_state_[2]\\\, B => 
        \Z\\SDram_rd_0_rd_state_[1]\\\, Y => N_383);
    
    \cs_n_1_RNO_1[0]\ : OR2A
      port map(A => \Z\\SDRAM_wr_0_wr_state_[2]\\\, B => N_370, Y
         => N_357);
    
    temp_w_n3_0_i_0 : XA1A
      port map(A => N_217, B => \temp_w[3]_net_1\, C => N_191, Y
         => \temp_w_n3_0_i_0\);
    
    \SD_wrAddr_row_RNO[0]\ : XA1A
      port map(A => N_7, B => \SD_wrAddr_row[0]_net_1\, C => 
        un7_sdram_enreg, Y => \SD_wrAddr_row_6[0]\);
    
    \SD_WrAddr_col[10]\ : DFN1E1C0
      port map(D => N_21, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => SD_WrAddr_cole, Q => 
        \SD_WrAddr_col[10]_net_1\);
    
    rdrow_end_RNO : NOR3C
      port map(A => un4lt10_i_a2_0_a7_2, B => un4lt10_i_a2_0_a7_1, 
        C => un4lt10_i_a2_0_a7_3, Y => N_565);
    
    dly1_SDoneFrameOk : DFN1C0
      port map(D => sd_wraddr_row20, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \dly1_SDoneFrameOk\);
    
    un1_SD_rdAddr_row_ADD_13x13_medium_area_I10_Y : OR3C
      port map(A => \SD_rdAddr_col[10]_net_1\, B => 
        \SD_rdAddr_row[0]_net_1\, C => \SD_rdAddr_row[1]_net_1\, 
        Y => N215);
    
    \SD_wrAddr_row_RNO[1]\ : XA1
      port map(A => \SD_wrAddr_row[1]_net_1\, B => N153, C => 
        un7_sdram_enreg, Y => \SD_wrAddr_row_6[1]\);
    
    \addr_RNO_1[10]\ : OR3C
      port map(A => N_186_0, B => N_211, C => N_223, Y => N_365);
    
    we_n_4_0_0_o4 : NOR2A
      port map(A => \Z\\Sdram_ini_0_ini_state_[0]\\\, B => 
        \Z\\Sdram_ini_0_ini_state_[1]\\\, Y => N_198);
    
    un1_SD_rdAddr_row_ADD_13x13_medium_area_I22_un1_Y_0 : NOR2B
      port map(A => \SD_rdAddr_row[11]_net_1\, B => N242_0, Y => 
        ADD_13x13_medium_area_I22_un1_Y_0);
    
    \SD_WrAddr_col_RNO[9]\ : XA1B
      port map(A => N_209, B => \SD_WrAddr_col[9]_net_1\, C => 
        un1_sdram_enreg_2, Y => N_19);
    
    \SD_WrAddr_col_RNI47BB[4]\ : OR3
      port map(A => \SD_WrAddr_col[3]_net_1\, B => 
        \SD_WrAddr_col[4]_net_1\, C => \SD_WrAddr_col[9]_net_1\, 
        Y => N_239);
    
    \SD_WrAddr_col_RNI7MI7[7]\ : OR2
      port map(A => \SD_WrAddr_col[7]_net_1\, B => 
        \SD_WrAddr_col[8]_net_1\, Y => 
        \un1_sd_wraddr_row8_i_o7_1[12]\);
    
    \SD_rdAddr_row_RNO[10]\ : XA1C
      port map(A => N199, B => N247, C => N_202, Y => 
        \SD_rdAddr_row_6[10]\);
    
    SDoneFrameOk : DFN1C0
      port map(D => \dly3_SDoneFrameOk\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => Sdram_cmd_0_SDoneFrameOk);
    
    un1_SD_wrAddr_row_ADD_13x13_medium_area_I22_un1_Y_1 : NOR3C
      port map(A => \SD_wrAddr_row[10]_net_1\, B => 
        \SD_wrAddr_row[11]_net_1\, C => N242, Y => 
        ADD_13x13_medium_area_I22_un1_Y_1);
    
    cas_n_RNO_0 : OR2
      port map(A => \Z\\Sdram_ini_0_ini_state_[1]\\\, B => 
        \Z\\Sdram_ini_0_ini_state_[2]\\\, Y => cas_n_4_6_0_a7_1_0);
    
    we_n : DFN1P0
      port map(D => we_n_4, CLK => PLL_Test1_0_Sys_66M_Clk, PRE
         => PLL_Test1_0_SysRst_O, Q => SD_we_n_c);
    
    \SD_WrAddr_col_RNO[7]\ : XA1B
      port map(A => N_199, B => \SD_WrAddr_col[7]_net_1\, C => 
        un1_sdram_enreg_2, Y => N_15);
    
    \SD_WrAddr_col_RNI92RL[10]\ : NOR2B
      port map(A => \SD_WrAddr_col[10]_net_1\, B => N_238, Y => 
        \un1_sd_wraddr_row8_i_0[12]\);
    
    \SD_rdAddr_row_RNI7CI7[12]\ : NOR3A
      port map(A => \SD_rdAddr_row[10]_net_1\, B => 
        \SD_rdAddr_row[12]_net_1\, C => \SD_rdAddr_row[8]_net_1\, 
        Y => sd_rdaddr_row18_0_a7_6);
    
    \SD_rdAddr_row[0]\ : DFN1C0
      port map(D => \SD_rdAddr_row_6[0]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \SD_rdAddr_row[0]_net_1\);
    
    \addr_RNO_3[10]\ : NOR3C
      port map(A => N_367, B => \addr_RNO_7[10]_net_1\, C => 
        N_364, Y => \addr_14_i_0_1[10]\);
    
    WFifo_re_RNO_1 : OR2
      port map(A => \temp_w[3]_net_1\, B => 
        \Z\\SDRAM_wr_0_wr_state_[1]\\\, Y => un1_cs_n7_4_i_0_a7_0);
    
    \SD_wrAddr_row[2]\ : DFN1C0
      port map(D => \SD_wrAddr_row_6[2]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \SD_wrAddr_row[2]_net_1\);
    
    \addr_RNO_5[7]\ : OR3A
      port map(A => N_186_0, B => N_192, C => 
        \SD_rdAddr_row[7]_net_1\, Y => N_331);
    
    \addr_RNO_5[5]\ : OR3B
      port map(A => N_186, B => \SD_rdAddr_row[5]_net_1\, C => 
        N_192, Y => N_320);
    
    un1_SD_wrAddr_row_ADD_13x13_medium_area_I35_un1_Y : OR2B
      port map(A => N258_0, B => \SD_wrAddr_row[6]_net_1\, Y => 
        I35_un1_Y_0);
    
    \SD_rdAddr_row_RNO[2]\ : XA1C
      port map(A => \SD_rdAddr_row[2]_net_1\, B => N215, C => 
        N_202, Y => \SD_rdAddr_row_6[2]\);
    
    \addr_RNO_7[10]\ : OR3A
      port map(A => \Z\\SDRAM_wr_0_wr_state_[0]\\\, B => 
        \Z\\SDRAM_wr_0_wr_state_[1]\\\, C => N_225, Y => 
        \addr_RNO_7[10]_net_1\);
    
    \SD_rdAddr_row[9]\ : DFN1C0
      port map(D => \SD_rdAddr_row_6[9]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \SD_rdAddr_row[9]_net_1\);
    
    ras_n_5_7_0_0_o4 : OR2A
      port map(A => \Z\\SDRAM_Ref_0_Ref_state_[0]\\\, B => 
        \Z\\SDRAM_Ref_0_Ref_state_[2]\\\, Y => N_187);
    
    \addr_RNO_2[0]\ : OR3B
      port map(A => N_186, B => \SD_addr_c[0]\, C => N_189, Y => 
        N_300);
    
    \SD_rdAddr_row[8]\ : DFN1C0
      port map(D => \SD_rdAddr_row_6[8]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \SD_rdAddr_row[8]_net_1\);
    
    un1_SD_wrAddr_row_ADD_13x13_medium_area_I22_Y : AO1
      port map(A => ADD_13x13_medium_area_I22_un1_Y_1, B => 
        N245_0, C => sd_wraddr_row20, Y => N237_0);
    
    \addr_RNO_0[8]\ : NOR3C
      port map(A => \addr_RNO_2[8]_net_1\, B => N_338, C => 
        \addr_RNO_4[8]_net_1\, Y => \addr_11_0_i_2[8]\);
    
    un1_SD_wrAddr_row_ADD_13x13_medium_area_I0_CO1 : NOR2A
      port map(A => \SD_wrAddr_row[0]_net_1\, B => N_7, Y => N153);
    
    \addr_RNO_1[4]\ : OA1
      port map(A => N_191, B => \SD_wrAddr_row[4]_net_1\, C => 
        \addr_RNO_5[4]_net_1\, Y => \addr_11_0_i_1[4]\);
    
    un1_SD_wrAddr_row_ADD_13x13_medium_area_I15_Y_1 : NOR3C
      port map(A => \SD_wrAddr_row[6]_net_1\, B => 
        \SD_wrAddr_row[7]_net_1\, C => N253, Y => 
        ADD_13x13_medium_area_I15_Y_1);
    
    \SD_wrAddr_row[9]\ : DFN1C0
      port map(D => \SD_wrAddr_row_6[9]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \SD_wrAddr_row[9]_net_1\);
    
    \addr_RNO_1[2]\ : OA1A
      port map(A => N_186_0, B => N_371, C => 
        \addr_RNO_4[2]_net_1\, Y => \addr_11_0_i_2[2]\);
    
    \SD_wrAddr_row_RNO[11]\ : XA1A
      port map(A => N261_i, B => ADD_13x13_medium_area_I48_Y_0_0, 
        C => un7_sdram_enreg, Y => \SD_wrAddr_row_6[11]\);
    
    sdram_enReg_RNI9B9H1 : OR3C
      port map(A => un7_sdram_enreg, B => N_261, C => N_372, Y
         => SD_WrAddr_cole);
    
    un1_SD_wrAddr_row_ADD_13x13_medium_area_I33_Y : AOI1
      port map(A => N247_0, B => \SD_wrAddr_row[10]_net_1\, C => 
        sd_wraddr_row20, Y => N261_i);
    
    \addr_RNO_3[2]\ : OR2
      port map(A => \SD_wrAddr_row[2]_net_1\, B => N_186, Y => 
        N_308);
    
    \addr_RNO_4[7]\ : OR3A
      port map(A => N_186_0, B => N_371, C => 
        \SD_rdAddr_col[7]_net_1\, Y => \addr_RNO_4[7]_net_1\);
    
    \addr_RNO_1[8]\ : OA1
      port map(A => N_191, B => \SD_wrAddr_row[8]_net_1\, C => 
        N_336, Y => \addr_11_0_i_1[8]\);
    
    \addr_RNO_0[12]\ : AOI1
      port map(A => N_384, B => \SD_addr_c[12]\, C => N_343_1, Y
         => N_343);
    
    un1_SD_rdAddr_row_ADD_13x13_medium_area_I49_Y_0_0 : XOR2
      port map(A => \SD_rdAddr_row[12]_net_1\, B => 
        sd_rdaddr_row18_i, Y => ADD_13x13_medium_area_I49_Y_0_0_0);
    
    \SD_rdAddr_row_RNIJS44[9]\ : NOR2
      port map(A => \SD_rdAddr_row[9]_net_1\, B => 
        \SD_rdAddr_row[11]_net_1\, Y => sd_rdaddr_row18_0_a7_4);
    
    un1_SD_wrAddr_row_ADD_13x13_medium_area_I8_Y : NOR2B
      port map(A => \SD_wrAddr_row[5]_net_1\, B => 
        \SD_wrAddr_row[4]_net_1\, Y => N253);
    
    \addr_RNO_3[5]\ : OR2A
      port map(A => \SD_WrAddr_col[5]_net_1\, B => N_372, Y => 
        N_323);
    
    \addr_RNO[12]\ : NOR3
      port map(A => N_343, B => N_345, C => N_344, Y => N_178);
    
    \addr[0]\ : DFN1C0
      port map(D => \addr_11[0]\, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \SD_addr_c[0]\);
    
    \dqm_4_iv_i_0_a7_0[0]\ : NOR3A
      port map(A => \Z\\SDRAM_wr_0_wr_state_[2]\\\, B => 
        \Z\\SDRAM_wr_0_wr_state_[0]\\\, C => 
        \Z\\SDRAM_wr_0_wr_state_[1]\\\, Y => N_264);
    
    \SD_WrAddr_col_RNO[4]\ : XA1B
      port map(A => \SD_WrAddr_col[3]_net_1\, B => 
        \SD_WrAddr_col[4]_net_1\, C => un1_sdram_enreg_2, Y => 
        N_9_i_0);
    
    \SD_rdAddr_col_RNO[5]\ : XA1B
      port map(A => N_195, B => \SD_rdAddr_col[5]_net_1\, C => 
        N_428, Y => N_35);
    
    \addr_RNO_1[9]\ : OA1
      port map(A => N_191, B => \SD_wrAddr_row[9]_net_1\, C => 
        N_251, Y => \addr_11_i_0_1[9]\);
    
    un1_SD_rdAddr_row_ADD_13x13_medium_area_I22_un1_Y_1 : NOR2B
      port map(A => ADD_13x13_medium_area_I22_un1_Y_0, B => N199, 
        Y => ADD_13x13_medium_area_I22_un1_Y_1_0);
    
    \addr_RNO_1[6]\ : OA1
      port map(A => N_191, B => \SD_wrAddr_row[6]_net_1\, C => 
        \addr_RNO_5[6]_net_1\, Y => \addr_11_0_i_1[6]\);
    
    \addr_RNO_1[5]\ : OA1A
      port map(A => \SD_wrAddr_row[5]_net_1\, B => N_191, C => 
        N_320, Y => \addr_11_i_i_1[5]\);
    
    un1_SD_wrAddr_row_ADD_13x13_medium_area_I48_Y_0_0 : XOR2
      port map(A => \SD_wrAddr_row[11]_net_1\, B => 
        sd_wraddr_row20, Y => ADD_13x13_medium_area_I48_Y_0_0);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \SD_WrAddr_col[7]\ : DFN1E1C0
      port map(D => N_15, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => SD_WrAddr_cole, Q => 
        \SD_WrAddr_col[7]_net_1\);
    
    \SD_rdAddr_row_RNO[11]\ : XA1C
      port map(A => N261, B => ADD_13x13_medium_area_I48_Y_0_0_0, 
        C => N_202, Y => \SD_rdAddr_row_6[11]\);
    
    \addr_RNO[8]\ : NOR3C
      port map(A => \addr_11_0_i_2[8]\, B => \addr_11_0_i_1[8]\, 
        C => N_249_i, Y => N_174_i_0);
    
    \addr[8]\ : DFN1C0
      port map(D => N_174_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \SD_addr_c[8]\);
    
    \SD_wrAddr_row[12]\ : DFN1C0
      port map(D => \SD_wrAddr_row_6[12]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \SD_wrAddr_row[12]_net_1\);
    
    \SD_WrAddr_col[4]\ : DFN1E1C0
      port map(D => N_9_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => SD_WrAddr_cole, Q => 
        \SD_WrAddr_col[4]_net_1\);
    
    \SD_rdAddr_col_RNO_0[10]\ : OR2B
      port map(A => \SD_rdAddr_col[9]_net_1\, B => N_214, Y => 
        N_219);
    
    we_n_RNO_4 : OR2A
      port map(A => N_189, B => N_370, Y => N_360);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    \SD_WrAddr_col_RNO[8]\ : XA1B
      port map(A => N_203, B => \SD_WrAddr_col[8]_net_1\, C => 
        un1_sdram_enreg_2, Y => N_17);
    
    \LVDS_enReg\ : DFN1C0
      port map(D => CMOS_DrvX_0_SDramEn, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => LVDS_enReg);
    
    \dqm_4_iv_i_0_a4[0]\ : OR2A
      port map(A => \Z\\SDRAM_wr_0_wr_state_[1]\\\, B => N_186_0, 
        Y => N_372);
    
    \SD_WrAddr_col_RNIE3GQ[9]\ : OR2B
      port map(A => \SD_WrAddr_col[9]_net_1\, B => N_209, Y => 
        N_218);
    
    \cs_n_1_RNO_3[0]\ : OR3C
      port map(A => N_187, B => \Z\\SDRAM_wr_0_wr_state_[1]\\\, C
         => N_186_0, Y => N_358);
    
    \SD_WrAddr_col[6]\ : DFN1E1C0
      port map(D => N_13, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => SD_WrAddr_cole, Q => 
        \SD_WrAddr_col[6]_net_1\);
    
    \SD_WrAddr_col[5]\ : DFN1E1C0
      port map(D => N_11_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => SD_WrAddr_cole, Q => 
        \SD_WrAddr_col[5]_net_1\);
    
    \dqm_1[0]\ : DFN1P0
      port map(D => \dqm_1_RNO[0]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, PRE => PLL_Test1_0_SysRst_O, Q
         => SD_dqm_c_c_c_c_c_c_c_c(1));
    
    \SD_rdAddr_row[10]\ : DFN1C0
      port map(D => \SD_rdAddr_row_6[10]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \SD_rdAddr_row[10]_net_1\);
    
    \SD_WrAddr_col[3]\ : DFN1E1C0
      port map(D => N_16, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => SD_WrAddr_cole, Q => 
        \SD_WrAddr_col[3]_net_1\);
    
    \addr_RNO_2[8]\ : OR3A
      port map(A => N_186_0, B => N_189, C => \SD_addr_c[8]\, Y
         => \addr_RNO_2[8]_net_1\);
    
    \SD_WrAddr_col[9]\ : DFN1E1C0
      port map(D => N_19, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => SD_WrAddr_cole, Q => 
        \SD_WrAddr_col[9]_net_1\);
    
    \addr_RNO_2[3]\ : OR3A
      port map(A => N_186, B => N_192, C => 
        \SD_rdAddr_row[3]_net_1\, Y => \addr_RNO_2[3]_net_1\);
    
    cas_n_RNO_5 : MX2
      port map(A => \Z\\SDRAM_wr_0_wr_state_[0]\\\, B => 
        \Z\\SDRAM_wr_0_wr_state_[2]\\\, S => 
        \Z\\SDRAM_wr_0_wr_state_[1]\\\, Y => N_231);
    
    \addr_RNO_2[12]\ : NOR3A
      port map(A => N_191, B => N_192, C => 
        \SD_rdAddr_row[12]_net_1\, Y => N_344);
    
    un1_SD_wrAddr_row_ADD_13x13_medium_area_I14_Y : NOR2B
      port map(A => ADD_13x13_medium_area_I14_Y_0, B => N215_0, Y
         => N256_0);
    
    \SD_rdAddr_row[5]\ : DFN1C0
      port map(D => \SD_rdAddr_row_6[5]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \SD_rdAddr_row[5]_net_1\);
    
    WFifo_re_RNO : OAI1
      port map(A => N_217, B => un1_cs_n7_4_i_0_a7_1, C => N_191, 
        Y => N_10);
    
    \SD_wrAddr_row[6]\ : DFN1C0
      port map(D => \SD_wrAddr_row_6[6]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \SD_wrAddr_row[6]_net_1\);
    
    \SD_rdAddr_row_RNIFTC1[3]\ : NOR2
      port map(A => \SD_rdAddr_row[2]_net_1\, B => 
        \SD_rdAddr_row[3]_net_1\, Y => sd_rdaddr_row18_0_a7_2);
    
    wrrow_end_RNO : OAI1
      port map(A => N_218, B => \SD_WrAddr_col[10]_net_1\, C => 
        N_248, Y => N_4);
    
    \SD_wrAddr_row[7]\ : DFN1C0
      port map(D => \SD_wrAddr_row_6[7]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \SD_wrAddr_row[7]_net_1\);
    
    \SD_WrAddr_col_RNO_0[5]\ : AO1
      port map(A => \SD_WrAddr_col[4]_net_1\, B => 
        \SD_WrAddr_col[3]_net_1\, C => \SD_WrAddr_col[5]_net_1\, 
        Y => N_255);
    
    \SD_rdAddr_col_RNIQLR61[7]\ : NOR3C
      port map(A => N_197, B => \SD_rdAddr_col[6]_net_1\, C => 
        \SD_rdAddr_col[7]_net_1\, Y => N_204);
    
    \addr_RNO_0[2]\ : AOI1B
      port map(A => \addr_11_0_i_a7_0[2]\, B => N_192, C => N_308, 
        Y => \addr_11_0_i_0[2]\);
    
    un1_SD_rdAddr_row_ADD_13x13_medium_area_I27_Y : OR2B
      port map(A => N245, B => N242_0, Y => N247);
    
    temp_w_n1_0_i_0 : XA1
      port map(A => \temp_w[0]_net_1\, B => \temp_w[1]_net_1\, C
         => N_191, Y => \temp_w_n1_0_i_0\);
    
    \addr[5]\ : DFN1C0
      port map(D => N_168, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \SD_addr_c[5]\);
    
    \SD_rdAddr_row_RNI9MI5[5]\ : NOR3A
      port map(A => sd_rdaddr_row18_0_a7_4, B => 
        \SD_rdAddr_row[7]_net_1\, C => \SD_rdAddr_row[5]_net_1\, 
        Y => sd_rdaddr_row18_0_a7_8);
    
    \addr_RNO_2[7]\ : OR3A
      port map(A => N_186_0, B => N_189, C => \SD_addr_c[7]\, Y
         => \addr_RNO_2[7]_net_1\);
    
    \addr_RNO[0]\ : OR3C
      port map(A => \addr_11_0_0_0[0]\, B => N_630, C => N_249_i, 
        Y => \addr_11[0]\);
    
    rdrow_end_RNO_1 : NOR2
      port map(A => \SD_rdAddr_col[6]_net_1\, B => 
        \SD_rdAddr_col[7]_net_1\, Y => un4lt10_i_a2_0_a7_1);
    
    un1_SD_wrAddr_row_ADD_13x13_medium_area_I36_un1_Y : OR2B
      port map(A => N256_0, B => \SD_wrAddr_row[4]_net_1\, Y => 
        I36_un1_Y_0);
    
    \SD_rdAddr_row_RNO[12]\ : XA1C
      port map(A => N237, B => ADD_13x13_medium_area_I49_Y_0_0_0, 
        C => N_202, Y => \SD_rdAddr_row_6[12]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \addr_RNO_4[9]\ : OR3A
      port map(A => N_186_0, B => N_371, C => 
        \SD_rdAddr_col[9]_net_1\, Y => \addr_RNO_4[9]_net_1\);
    
    \addr[1]\ : DFN1C0
      port map(D => \addr_11[1]\, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \SD_addr_c[1]\);
    
    \SD_rdAddr_col_RNO[10]\ : NOR3
      port map(A => N_219, B => N_428, C => N_371, Y => 
        \SD_rdAddr_col_RNO[10]_net_1\);
    
    \SD_rdAddr_col_RNI13HF[3]\ : NOR2B
      port map(A => \SD_rdAddr_col[4]_net_1\, B => 
        \SD_rdAddr_col[3]_net_1\, Y => N_195);
    
    \SD_wrAddr_row[10]\ : DFN1C0
      port map(D => \SD_wrAddr_row_6[10]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \SD_wrAddr_row[10]_net_1\);
    
    WFifo_re : DFN1E1C0
      port map(D => \Z\\SDRAM_wr_0_wr_state_[0]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => N_10, Q => Sdram_cmd_0_WFifo_re);
    
    un1_SD_rdAddr_row_ADD_13x13_medium_area_I6_Y : NOR2B
      port map(A => \SD_rdAddr_row[9]_net_1\, B => 
        \SD_rdAddr_row[8]_net_1\, Y => N242_0);
    
    ras_n_RNO_1 : AOI1B
      port map(A => N_221, B => N_187, C => N_635, Y => 
        ras_n_5_7_0_0_0);
    
    \addr_RNO_1[11]\ : NOR2
      port map(A => \SD_wrAddr_row[11]_net_1\, B => N_191, Y => 
        N_342);
    
    \addr_RNO_0[6]\ : NOR3C
      port map(A => \addr_RNO_2[6]_net_1\, B => 
        \addr_RNO_3[6]_net_1\, C => \addr_RNO_4[6]_net_1\, Y => 
        \addr_11_0_i_2[6]\);
    
    un1_SD_rdAddr_row_ADD_13x13_medium_area_I14_Y : NOR2
      port map(A => ADD_13x13_medium_area_I14_Y_0_0, B => N215, Y
         => N256);
    
    \SD_WrAddr_col_RNO[3]\ : NOR2
      port map(A => un1_sdram_enreg_2, B => 
        \SD_WrAddr_col[3]_net_1\, Y => N_16);
    
    \addr_RNO_5[3]\ : OR2
      port map(A => \SD_wrAddr_row[3]_net_1\, B => N_191, Y => 
        \addr_RNO_5[3]_net_1\);
    
    \addr_RNO_2[6]\ : OR3A
      port map(A => N_186, B => N_189, C => \SD_addr_c[6]\, Y => 
        \addr_RNO_2[6]_net_1\);
    
    \SD_wrAddr_row[1]\ : DFN1C0
      port map(D => \SD_wrAddr_row_6[1]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \SD_wrAddr_row[1]_net_1\);
    
    \SD_wrAddr_row_RNIT9BC[2]\ : NOR2A
      port map(A => \SD_wrAddr_row[10]_net_1\, B => 
        \SD_wrAddr_row[2]_net_1\, Y => sd_wraddr_row20_0_a7_4);
    
    \addr_RNO_0[5]\ : NOR3C
      port map(A => N_319, B => N_323, C => N_322, Y => 
        \addr_11_i_i_2[5]\);
    
    \SD_rdAddr_row_RNIUUBH[1]\ : OR3C
      port map(A => sd_rdaddr_row18_0_a7_8, B => 
        sd_rdaddr_row18_0_a7_7, C => sd_rdaddr_row18_0_a7_9, Y
         => sd_rdaddr_row18_i);
    
    \temp_w[2]\ : DFN1C0
      port map(D => \temp_w_n2_0_i_0\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \temp_w[2]_net_1\);
    
    we_n_RNO_0 : NOR3C
      port map(A => \we_n_RNO_2\, B => N_362, C => N_360, Y => 
        we_n_4_0_0_1);
    
    un1_SD_rdAddr_row_ADD_13x13_medium_area_I33_Y : AO1C
      port map(A => N247, B => \SD_rdAddr_row[10]_net_1\, C => 
        sd_rdaddr_row18_i, Y => N261);
    
    \SD_rdAddr_col_RNO[6]\ : XA1B
      port map(A => N_197, B => \SD_rdAddr_col[6]_net_1\, C => 
        N_428, Y => N_541);
    
    \temp_w[3]\ : DFN1C0
      port map(D => \temp_w_n3_0_i_0\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \temp_w[3]_net_1\);
    
    cas_n_RNO_2 : OR3A
      port map(A => \Z\\SDram_rd_0_rd_state_[1]\\\, B => N_220, C
         => N_370, Y => N_637);
    
    dly3_SDoneFrameOk : DFN1C0
      port map(D => \dly2_SDoneFrameOk\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \dly3_SDoneFrameOk\);
    
    un1_SD_wrAddr_row_ADD_13x13_medium_area_I6_Y : NOR2B
      port map(A => \SD_wrAddr_row[9]_net_1\, B => 
        \SD_wrAddr_row[8]_net_1\, Y => N242);
    
    cas_n_RNO_4 : OR3A
      port map(A => N_193, B => N_201, C => N_370, Y => N_638);
    
    we_n_RNO : OR3C
      port map(A => N_216, B => we_n_4_0_0_1, C => N_361, Y => 
        we_n_4);
    
    un1_SD_wrAddr_row_ADD_13x13_medium_area_I47_Y_0_0 : XOR2
      port map(A => \SD_wrAddr_row[10]_net_1\, B => 
        sd_wraddr_row20, Y => ADD_13x13_medium_area_I47_Y_0_0);
    
    cas_n_4_6_0_0_o4 : OR2A
      port map(A => \Z\\SDram_rd_0_rd_state_[2]\\\, B => 
        \Z\\SDram_rd_0_rd_state_[0]\\\, Y => N_193);
    
    \dqm_4_iv_i_0_a7_0_2[0]\ : NOR3A
      port map(A => \Z\\SDRAM_wr_0_wr_state_[2]\\\, B => 
        \Z\\SDRAM_wr_0_wr_state_[0]\\\, C => 
        \Z\\SDRAM_wr_0_wr_state_[1]\\\, Y => N_264_2);
    
    \SD_wrAddr_row_RNO[10]\ : XA1
      port map(A => N247_0, B => ADD_13x13_medium_area_I47_Y_0_0, 
        C => un7_sdram_enreg, Y => \SD_wrAddr_row_6[10]\);
    
    ras_n_5_7_0_0_a2 : OR2A
      port map(A => N_187, B => \Z\\SDRAM_wr_0_wr_state_[0]\\\, Y
         => N_370);
    
    \SD_rdAddr_row_RNO[8]\ : XA1B
      port map(A => \SD_rdAddr_row[8]_net_1\, B => N245, C => 
        N_202, Y => \SD_rdAddr_row_6[8]\);
    
    \SD_rdAddr_col_RNO[9]\ : XA1B
      port map(A => N_214, B => \SD_rdAddr_col[9]_net_1\, C => 
        N_428, Y => N_544);
    
    \SD_wrAddr_row_RNO[4]\ : XA1
      port map(A => \SD_wrAddr_row[4]_net_1\, B => N256_0, C => 
        un7_sdram_enreg, Y => \SD_wrAddr_row_6[4]\);
    
    \SD_rdAddr_col_RNO[4]\ : XA1B
      port map(A => \SD_rdAddr_col[3]_net_1\, B => 
        \SD_rdAddr_col[4]_net_1\, C => N_428, Y => N_540);
    
    \SD_WrAddr_col_RNI36I7[5]\ : OR2
      port map(A => \SD_WrAddr_col[5]_net_1\, B => 
        \SD_WrAddr_col[6]_net_1\, Y => 
        \un1_sd_wraddr_row8_i_o7_0[12]\);
    
    \SD_rdAddr_col_RNO[7]\ : NOR3
      port map(A => N_204, B => N_297, C => N_428, Y => N_542);
    
    \addr[9]\ : DFN1C0
      port map(D => N_6_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \SD_addr_c[9]\);
    
    we_n_RNO_1 : OR2A
      port map(A => N_187, B => N_191, Y => N_361);
    
    \SD_WrAddr_col_RNID9611[10]\ : OR2A
      port map(A => \un1_sd_wraddr_row8_i_0[12]\, B => N_239, Y
         => N_261);
    
    \cs_n_1_RNO_4[0]\ : XO1A
      port map(A => \Z\\SDRAM_Ref_0_Ref_state_[1]\\\, B => 
        \Z\\SDRAM_Ref_0_Ref_state_[2]\\\, C => 
        \Z\\SDRAM_Ref_0_Ref_state_[0]\\\, Y => 
        \cs_n_1_RNO_4[0]_net_1\);
    
    \addr_RNO[6]\ : NOR3C
      port map(A => \addr_11_0_i_2[6]\, B => \addr_11_0_i_1[6]\, 
        C => N_249_i, Y => N_170_i_0);
    
    un1_SD_rdAddr_row_ADD_13x13_medium_area_I38_Y_0 : AX1E
      port map(A => \SD_rdAddr_col[10]_net_1\, B => 
        \SD_rdAddr_row[0]_net_1\, C => \SD_rdAddr_row[1]_net_1\, 
        Y => \un1_SD_rdAddr_row_i[1]\);
    
    un1_SD_wrAddr_row_ADD_13x13_medium_area_I27_Y : NOR2B
      port map(A => N245_0, B => N242, Y => N247_0);
    
    \SD_rdAddr_row_RNO[1]\ : NOR2
      port map(A => \un1_SD_rdAddr_row_i[1]\, B => N_202, Y => 
        \SD_rdAddr_row_6[1]\);
    
    SD_rdAddr_collde_0_0_a4 : OR2
      port map(A => N_193, B => \Z\\SDram_rd_0_rd_state_[1]\\\, Y
         => N_371);
    
    \addr_11_0_i_o4[2]\ : OR2A
      port map(A => \Z\\SDRAM_wr_0_wr_state_[0]\\\, B => 
        \Z\\SDRAM_wr_0_wr_state_[2]\\\, Y => N_186);
    
    \addr_RNO_5[8]\ : OR3A
      port map(A => N_186_0, B => N_192, C => 
        \SD_rdAddr_row[8]_net_1\, Y => N_336);
    
    \SD_WrAddr_col_RNO[10]\ : XA1C
      port map(A => N_218, B => \SD_WrAddr_col[10]_net_1\, C => 
        un1_sdram_enreg_2, Y => N_21);
    
    \addr_RNO_2[2]\ : AOI1B
      port map(A => N_384, B => \SD_addr_c[2]\, C => N_186_0, Y
         => \addr_11_0_i_a7_0[2]\);
    
    \SD_rdAddr_col[8]\ : DFN1E1C0
      port map(D => N_543, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => SD_rdAddr_cole, Q => 
        \SD_rdAddr_col[8]_net_1\);
    
    \addr_RNO_8[10]\ : OR3B
      port map(A => N_224, B => N_186_0, C => N_193, Y => N_364);
    
    \SD_wrAddr_row_RNI9H2H[12]\ : NOR3
      port map(A => \SD_wrAddr_row[0]_net_1\, B => 
        \SD_wrAddr_row[12]_net_1\, C => \SD_wrAddr_row[8]_net_1\, 
        Y => sd_wraddr_row20_0_a7_6);
    
    ras_n_RNO_0 : OR3A
      port map(A => N_190, B => N_201, C => N_370, Y => N_634);
    
    \addr_RNO[7]\ : NOR3C
      port map(A => \addr_11_0_i_2[7]\, B => \addr_11_0_i_1[7]\, 
        C => N_249_i, Y => N_172_i_0);
    
    \SD_rdAddr_row_RNO[0]\ : XA1C
      port map(A => N_539, B => \SD_rdAddr_row[0]_net_1\, C => 
        N_202, Y => \SD_rdAddr_row_6[0]\);
    
    temp_w_n0_0_i_0 : NOR2A
      port map(A => N_191, B => \temp_w[0]_net_1\, Y => 
        \temp_w_n0_0_i_0\);
    
    \addr_RNO_4[3]\ : OA1
      port map(A => N_372, B => \SD_WrAddr_col[3]_net_1\, C => 
        \addr_RNO_5[3]_net_1\, Y => \addr_11_0_i_0[3]\);
    
    \addr_RNO_5[6]\ : OR3A
      port map(A => N_186, B => N_192, C => 
        \SD_rdAddr_row[6]_net_1\, Y => \addr_RNO_5[6]_net_1\);
    
    \SD_rdAddr_row_RNO[3]\ : XA1B
      port map(A => \SD_rdAddr_row[3]_net_1\, B => I37_un1_Y, C
         => N_202, Y => \SD_rdAddr_row_6[3]\);
    
    \SD_WrAddr_col_RNIAS4F[5]\ : NOR2
      port map(A => \un1_sd_wraddr_row8_i_o7_1[12]\, B => 
        \un1_sd_wraddr_row8_i_o7_0[12]\, Y => N_238);
    
    rdrow_end : DFN1E0C0
      port map(D => \SD_rdAddr_col[10]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => N_565, Q => Sdram_cmd_0_rdrow_end);
    
    \SD_WrAddr_col_RNI55TI[7]\ : NOR2B
      port map(A => \SD_WrAddr_col[7]_net_1\, B => N_199, Y => 
        N_203);
    
    ras_n_5_7_0_a4_0 : NOR3C
      port map(A => \Z\\SDRAM_wr_0_wr_state_[1]\\\, B => 
        \Z\\SDRAM_wr_0_wr_state_[2]\\\, C => N_187, Y => N_379);
    
    \addr_RNO_3[6]\ : OR2
      port map(A => \SD_WrAddr_col[6]_net_1\, B => N_372, Y => 
        \addr_RNO_3[6]_net_1\);
    
    \dqm_4_iv_i_0_o4[0]\ : NOR2B
      port map(A => \Z\\SDRAM_wr_0_wr_state_[1]\\\, B => 
        \Z\\SDRAM_wr_0_wr_state_[0]\\\, Y => N_221);
    
    \cs_n_1_RNO_2[0]\ : OR3
      port map(A => N_201, B => N_370, C => N_205, Y => N_356);
    
    \SD_wrAddr_row_RNO[9]\ : XA1A
      port map(A => \SD_wrAddr_row[9]_net_1\, B => I34_un1_Y, C
         => un7_sdram_enreg, Y => \SD_wrAddr_row_6[9]\);
    
    \dqm_4_iv_i_0_a7_0_1[0]\ : NOR3A
      port map(A => \Z\\SDRAM_wr_0_wr_state_[2]\\\, B => 
        \Z\\SDRAM_wr_0_wr_state_[0]\\\, C => 
        \Z\\SDRAM_wr_0_wr_state_[1]\\\, Y => N_264_1);
    
    ras_n_5_7_0_0_o7 : OA1B
      port map(A => N_353_2, B => N_383, C => N_379, Y => N_216);
    
    dly2_SDoneFrameOk : DFN1C0
      port map(D => \dly1_SDoneFrameOk\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \dly2_SDoneFrameOk\);
    
    \addr_RNO_4[10]\ : MX2A
      port map(A => \SD_addr_c[10]\, B => 
        \Z\\Sdram_ini_0_ini_state_[2]\\\, S => N_198, Y => N_211);
    
    sdram_enReg_RNI0TAC : OR2A
      port map(A => \sdram_enReg\, B => CMOS_DrvX_0_LVDSen_2, Y
         => un7_sdram_enreg);
    
    \addr_11_0_i_o4_0_0[2]\ : OR2A
      port map(A => \Z\\SDRAM_wr_0_wr_state_[0]\\\, B => 
        \Z\\SDRAM_wr_0_wr_state_[2]\\\, Y => N_186_0);
    
    \addr_RNO_1[12]\ : NOR2
      port map(A => \SD_wrAddr_row[12]_net_1\, B => N_191, Y => 
        N_345);
    
    \SD_WrAddr_col_RNI0NAB[5]\ : OR3C
      port map(A => \SD_WrAddr_col[3]_net_1\, B => 
        \SD_WrAddr_col[4]_net_1\, C => \SD_WrAddr_col[5]_net_1\, 
        Y => N_196);
    
    \addr_RNO_5[4]\ : OR3A
      port map(A => N_186, B => N_192, C => 
        \SD_rdAddr_row[4]_net_1\, Y => \addr_RNO_5[4]_net_1\);
    
    \SD_wrAddr_row_RNO[2]\ : XA1
      port map(A => \SD_wrAddr_row[2]_net_1\, B => N215_0, C => 
        un7_sdram_enreg, Y => \SD_wrAddr_row_6[2]\);
    
    \SD_wrAddr_row[11]\ : DFN1C0
      port map(D => \SD_wrAddr_row_6[11]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \SD_wrAddr_row[11]_net_1\);
    
    \SD_wrAddr_row[5]\ : DFN1C0
      port map(D => \SD_wrAddr_row_6[5]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \SD_wrAddr_row[5]_net_1\);
    
    \SD_rdAddr_col_RNO[8]\ : XA1B
      port map(A => N_204, B => \SD_rdAddr_col[8]_net_1\, C => 
        N_428, Y => N_543);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    \SD_rdAddr_row_RNO[9]\ : XA1C
      port map(A => \SD_rdAddr_row[9]_net_1\, B => I34_un1_Y_0, C
         => N_202, Y => \SD_rdAddr_row_6[9]\);
    
    cas_n : DFN1P0
      port map(D => cas_n_4, CLK => PLL_Test1_0_Sys_66M_Clk, PRE
         => PLL_Test1_0_SysRst_O, Q => SD_cas_n_c);
    
    \addr_RNO_5[9]\ : OR3A
      port map(A => N_186_0, B => N_192, C => 
        \SD_rdAddr_row[9]_net_1\, Y => N_251);
    
    un1_cs_n7_4_i_0_o4 : OR2
      port map(A => N_186_0, B => \Z\\SDRAM_wr_0_wr_state_[1]\\\, 
        Y => N_191);
    
    \addr_11_0_i_a7_1_0[12]\ : OR2B
      port map(A => N_192, B => N_191, Y => N_343_1);
    
    Rfifo_weEN : DFN1E1
      port map(D => un1_rfifo_ween2_3, CLK => 
        PLL_Test1_0_Sys_66M_Clk, E => PLL_Test1_0_SysRst_O, Q => 
        \Rfifo_weEN\);
    
    rdrow_end_RNO_0 : NOR2
      port map(A => \SD_rdAddr_col[8]_net_1\, B => 
        \SD_rdAddr_col[9]_net_1\, Y => un4lt10_i_a2_0_a7_2);
    
    \SD_rdAddr_col_RNIQBON[10]\ : OR2
      port map(A => \SD_rdAddr_col[10]_net_1\, B => N_202, Y => 
        N_428);
    
    \addr_RNO_0[10]\ : NOR3C
      port map(A => N_365, B => N_366, C => \addr_14_i_0_1[10]\, 
        Y => \addr_14_i_0_3[10]\);
    
    \addr_RNO_0[4]\ : NOR3C
      port map(A => \addr_RNO_2[4]_net_1\, B => 
        \addr_RNO_3[4]_net_1\, C => \addr_RNO_4[4]_net_1\, Y => 
        \addr_11_0_i_2[4]\);
    
    \SD_rdAddr_row_RNO[5]\ : XA1C
      port map(A => \SD_rdAddr_row[5]_net_1\, B => I36_un1_Y, C
         => N_202, Y => \SD_rdAddr_row_6[5]\);
    
    \SD_rdAddr_row_RNO[7]\ : XA1C
      port map(A => \SD_rdAddr_row[7]_net_1\, B => I35_un1_Y, C
         => N_202, Y => \SD_rdAddr_row_6[7]\);
    
    \SD_wrAddr_row[0]\ : DFN1C0
      port map(D => \SD_wrAddr_row_6[0]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \SD_wrAddr_row[0]_net_1\);
    
    \SD_wrAddr_row_RNIKEE9[5]\ : NOR2
      port map(A => \SD_wrAddr_row[5]_net_1\, B => 
        \SD_wrAddr_row[7]_net_1\, Y => sd_wraddr_row20_0_a7_2);
    
    sdram_enReg_RNID6HD1 : OR2B
      port map(A => un7_sdram_enreg, B => N_261, Y => 
        un1_sdram_enreg_2);
    
    \addr_RNO_6[10]\ : OR2
      port map(A => N_187, B => \Z\\SDRAM_Ref_0_Ref_state_[1]\\\, 
        Y => N_367);
    
    \addr_RNO[3]\ : NOR3C
      port map(A => \addr_11_0_i_2[3]\, B => 
        \addr_RNO_1[3]_net_1\, C => N_249_i, Y => N_164_i_0);
    
    un1_SD_rdAddr_row_ADD_13x13_medium_area_I34_un1_Y : OR2B
      port map(A => N245, B => \SD_rdAddr_row[8]_net_1\, Y => 
        I34_un1_Y_0);
    
    \SD_rdAddr_col_RNIJQ9N[5]\ : NOR2B
      port map(A => \SD_rdAddr_col[5]_net_1\, B => N_195, Y => 
        N_197);
    
    \addr_RNO_3[9]\ : OR2
      port map(A => \SD_WrAddr_col[9]_net_1\, B => N_372, Y => 
        N_253);
    
    \addr_RNO[4]\ : NOR3C
      port map(A => \addr_11_0_i_2[4]\, B => \addr_11_0_i_1[4]\, 
        C => N_249_i, Y => N_166_i_0);
    
    \SD_rdAddr_row_RNO[4]\ : XA1B
      port map(A => \SD_rdAddr_row[4]_net_1\, B => N256, C => 
        N_202, Y => \SD_rdAddr_row_6[4]\);
    
    \addr_RNO_2[1]\ : OR3B
      port map(A => N_186, B => \SD_addr_c[1]\, C => N_189, Y => 
        N_303);
    
    un1_SD_rdAddr_row_ADD_13x13_medium_area_I15_Y : NOR2B
      port map(A => ADD_13x13_medium_area_I15_Y_1_0, B => N256, Y
         => N245);
    
    \cs_n_1_RNO[0]\ : OR3C
      port map(A => \cs_n_5_0_iv_0_0_1[0]\, B => N_357, C => 
        N_356, Y => \cs_n_5[0]\);
    
    \addr_RNO_1[1]\ : OR3B
      port map(A => N_186_0, B => \SD_rdAddr_row[1]_net_1\, C => 
        N_192, Y => N_304);
    
    \addr_RNO_4[4]\ : OR3A
      port map(A => N_186, B => N_371, C => 
        \SD_rdAddr_col[4]_net_1\, Y => \addr_RNO_4[4]_net_1\);
    
    \addr_RNO_3[3]\ : OR3A
      port map(A => N_186, B => N_189, C => \SD_addr_c[3]\, Y => 
        \addr_RNO_3[3]_net_1\);
    
    temp_w_n1_0_i_0_o4 : NOR2B
      port map(A => \temp_w[1]_net_1\, B => \temp_w[0]_net_1\, Y
         => N_207);
    
    \SD_wrAddr_row_RNI2GNO[9]\ : NOR3A
      port map(A => sd_wraddr_row20_0_a7_4, B => 
        \SD_wrAddr_row[11]_net_1\, C => \SD_wrAddr_row[9]_net_1\, 
        Y => sd_wraddr_row20_0_a7_8);
    
    \addr[12]\ : DFN1C0
      port map(D => N_178, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \SD_addr_c[12]\);
    
    \SD_wrAddr_row[8]\ : DFN1C0
      port map(D => \SD_wrAddr_row_6[8]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \SD_wrAddr_row[8]_net_1\);
    
    un1_SD_rdAddr_row_ADD_13x13_medium_area_I1_S_0 : XNOR2
      port map(A => sd_rdaddr_row18_i, B => 
        \SD_rdAddr_row[10]_net_1\, Y => N199);
    
    \addr_RNO[9]\ : NOR3C
      port map(A => \addr_11_i_0_2[9]\, B => \addr_11_i_0_1[9]\, 
        C => N_249_i, Y => N_6_i_0);
    
    \addr[4]\ : DFN1C0
      port map(D => N_166_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \SD_addr_c[4]\);
    
    un1_SD_wrAddr_row_ADD_13x13_medium_area_I37_un1_Y : OR2B
      port map(A => N215_0, B => \SD_wrAddr_row[2]_net_1\, Y => 
        I37_un1_Y_0);
    
    \addr_RNO_3[4]\ : OR2
      port map(A => \SD_WrAddr_col[4]_net_1\, B => N_372, Y => 
        \addr_RNO_3[4]_net_1\);
    
    \SD_rdAddr_row[4]\ : DFN1C0
      port map(D => \SD_rdAddr_row_6[4]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \SD_rdAddr_row[4]_net_1\);
    
    \SD_rdAddr_row_RNO_0[0]\ : OR2B
      port map(A => sd_rdaddr_row18_i, B => 
        \SD_rdAddr_col[10]_net_1\, Y => N_539);
    
    wrrow_end_RNO_0 : OR3A
      port map(A => N_238, B => N_239, C => 
        \SD_WrAddr_col[10]_net_1\, Y => N_248);
    
    \addr_RNO_2[5]\ : OR3B
      port map(A => N_186, B => \SD_addr_c[5]\, C => N_189, Y => 
        N_319);
    
    \addr[2]\ : DFN1C0
      port map(D => N_162_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \SD_addr_c[2]\);
    
    un1_SD_rdAddr_row_ADD_13x13_medium_area_I8_Y : NOR2B
      port map(A => \SD_rdAddr_row[5]_net_1\, B => 
        \SD_rdAddr_row[4]_net_1\, Y => N253_0);
    
    temp_w_n2_0_i_0_o4 : OR2B
      port map(A => \temp_w[2]_net_1\, B => N_207, Y => N_217);
    
    un1_SD_rdAddr_row_ADD_13x13_medium_area_I48_Y_0_0 : XOR2
      port map(A => \SD_rdAddr_row[11]_net_1\, B => 
        sd_rdaddr_row18_i, Y => ADD_13x13_medium_area_I48_Y_0_0_0);
    
    \SD_rdAddr_col_RNIEA451[10]\ : OR2A
      port map(A => N_371, B => N_428, Y => SD_rdAddr_cole);
    
    \addr_RNO_2[10]\ : OR3A
      port map(A => N_186_0, B => N_190, C => 
        \SD_rdAddr_row[10]_net_1\, Y => N_366);
    
    UU : WaveGenSingleZ18
      port map(Sdram_cmd_0_RFifo_we => Sdram_cmd_0_RFifo_we, 
        PLL_Test1_0_SysRst_O => PLL_Test1_0_SysRst_O, 
        PLL_Test1_0_Sys_66M_Clk => PLL_Test1_0_Sys_66M_Clk, 
        Rfifo_weEN => \Rfifo_weEN\);
    
    \addr[10]\ : DFN1C0
      port map(D => N_12_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \SD_addr_c[10]\);
    
    \SD_rdAddr_col_RNO[3]\ : NOR2
      port map(A => \SD_rdAddr_col[3]_net_1\, B => N_428, Y => 
        SD_rdAddr_col_n0);
    
    un1_SD_wrAddr_row_ADD_13x13_medium_area_I34_un1_Y : OR2B
      port map(A => N245_0, B => \SD_wrAddr_row[8]_net_1\, Y => 
        I34_un1_Y);
    
    un1_SD_wrAddr_row_ADD_13x13_medium_area_I14_Y_0 : NOR2B
      port map(A => \SD_wrAddr_row[3]_net_1\, B => 
        \SD_wrAddr_row[2]_net_1\, Y => 
        ADD_13x13_medium_area_I14_Y_0);
    
    \SD_wrAddr_row_RNIT4462[1]\ : NOR3C
      port map(A => sd_wraddr_row20_0_a7_8, B => 
        sd_wraddr_row20_0_a7_7, C => sd_wraddr_row20_0_a7_9, Y
         => sd_wraddr_row20);
    
    ras_n_RNO_2 : OR2
      port map(A => N_371, B => N_370, Y => N_635);
    
    \addr_RNO_10[10]\ : OR2A
      port map(A => \SD_rdAddr_col[10]_net_1\, B => 
        \Z\\SDram_rd_0_rd_state_[1]\\\, Y => N_224);
    
    \SD_rdAddr_row_RNO[6]\ : XA1B
      port map(A => \SD_rdAddr_row[6]_net_1\, B => N258, C => 
        N_202, Y => \SD_rdAddr_row_6[6]\);
    
    \addr_11_0_i_o4_0[2]\ : OR2
      port map(A => N_190, B => \Z\\SDram_rd_0_rd_state_[2]\\\, Y
         => N_192);
    
    un1_SD_rdAddr_row_ADD_13x13_medium_area_I36_un1_Y : OR2B
      port map(A => N256, B => \SD_rdAddr_row[4]_net_1\, Y => 
        I36_un1_Y);
    
    \temp_w[0]\ : DFN1C0
      port map(D => \temp_w_n0_0_i_0\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \temp_w[0]_net_1\);
    
    \SD_rdAddr_row_RNIRTV8[4]\ : NOR3A
      port map(A => sd_rdaddr_row18_0_a7_6, B => 
        \SD_rdAddr_row[6]_net_1\, C => \SD_rdAddr_row[4]_net_1\, 
        Y => sd_rdaddr_row18_0_a7_9);
    
    \SD_rdAddr_row[11]\ : DFN1C0
      port map(D => \SD_rdAddr_row_6[11]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \SD_rdAddr_row[11]_net_1\);
    
    un1_SD_wrAddr_row_ADD_13x13_medium_area_I15_Y : NOR2B
      port map(A => ADD_13x13_medium_area_I15_Y_1, B => N256_0, Y
         => N245_0);
    
    cas_n_4_6_0_a7_1_2 : OR2A
      port map(A => N_193, B => N_370, Y => N_353_2);
    
    \addr_RNO[10]\ : OA1
      port map(A => N_372, B => \SD_WrAddr_col[10]_net_1\, C => 
        \addr_14_i_0_3[10]\, Y => N_12_i_0);
    
    we_n_RNO_2 : OR3A
      port map(A => N_190, B => N_198, C => N_370, Y => 
        \we_n_RNO_2\);
    
    \cs_n_1_RNO_5[0]\ : OR3B
      port map(A => N_205, B => \Z\\SDram_rd_0_rd_state_[0]\\\, C
         => N_370, Y => N_355);
    
    \addr_RNO_1[0]\ : OR3B
      port map(A => N_186, B => \SD_rdAddr_row[0]_net_1\, C => 
        N_192, Y => N_630);
    
    \SD_Clk_1[1]\ : NOR2B
      port map(A => SD_cke_c_c(0), B => PLL_Test1_0_Sdram_clk, Y
         => SD_Clk_c_c(1));
    
    \SD_WrAddr_col_RNIAEA73[10]\ : OR2A
      port map(A => \un1_sd_wraddr_row8_i_1[12]\, B => 
        sd_wraddr_row20, Y => N_7);
    
    \addr_RNO_0[7]\ : NOR3C
      port map(A => \addr_RNO_2[7]_net_1\, B => N_333, C => 
        \addr_RNO_4[7]_net_1\, Y => \addr_11_0_i_2[7]\);
    
    un1_SD_wrAddr_row_ADD_13x13_medium_area_I49_Y_0_0 : XOR2
      port map(A => \SD_wrAddr_row[12]_net_1\, B => 
        sd_wraddr_row20, Y => ADD_13x13_medium_area_I49_Y_0_0);
    
    \SD_wrAddr_row[3]\ : DFN1C0
      port map(D => \SD_wrAddr_row_6[3]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \SD_wrAddr_row[3]_net_1\);
    
    un1_SD_rdAddr_row_ADD_13x13_medium_area_I37_un1_Y : NOR2A
      port map(A => \SD_rdAddr_row[2]_net_1\, B => N215, Y => 
        I37_un1_Y);
    
    \SD_rdAddr_col_RNIFPKE1[8]\ : NOR2B
      port map(A => \SD_rdAddr_col[8]_net_1\, B => N_204, Y => 
        N_214);
    
    \addr_RNO_4[5]\ : OR3B
      port map(A => N_186, B => \SD_rdAddr_col[5]_net_1\, C => 
        N_371, Y => N_322);
    
    sdram_enReg : DFN1C0
      port map(D => CMOS_DrvX_0_LVDSen, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \sdram_enReg\);
    
    ras_n_5_7_0_0_o2 : AOI1B
      port map(A => \Z\\Sdram_ini_0_ini_state_[2]\\\, B => 
        \Z\\Sdram_ini_0_ini_state_[1]\\\, C => 
        \Z\\Sdram_ini_0_ini_state_[0]\\\, Y => N_201);
    
    un1_rfifo_ween2_3_0_0_o4 : OR2
      port map(A => \Z\\SDram_rd_0_rd_state_[2]\\\, B => 
        \Z\\SDram_rd_0_rd_state_[1]\\\, Y => N_205);
    
    \addr_RNO_5[10]\ : OR2A
      port map(A => N_205, B => \Z\\SDram_rd_0_rd_state_[0]\\\, Y
         => N_223);
    
    \SD_wrAddr_row_RNO[6]\ : XA1
      port map(A => \SD_wrAddr_row[6]_net_1\, B => N258_0, C => 
        un7_sdram_enreg, Y => \SD_wrAddr_row_6[6]\);
    
    \addr[6]\ : DFN1C0
      port map(D => N_170_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \SD_addr_c[6]\);
    
    un1_SD_rdAddr_row_ADD_13x13_medium_area_I35_un1_Y : OR2B
      port map(A => N258, B => \SD_rdAddr_row[6]_net_1\, Y => 
        I35_un1_Y);
    
    cas_n_RNO_3 : MX2B
      port map(A => \Z\\SDRAM_Ref_0_Ref_state_[1]\\\, B => N_231, 
        S => N_187, Y => N_241);
    
    we_n_4_0_0_o2 : NOR3B
      port map(A => N_383, B => N_205, C => 
        \Z\\SDram_rd_0_rd_state_[0]\\\, Y => N_189);
    
    un1_SD_rdAddr_row_ADD_13x13_medium_area_I32_Y : NOR2B
      port map(A => N256, B => N253_0, Y => N258);
    
    \SD_WrAddr_col[8]\ : DFN1E1C0
      port map(D => N_17, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => SD_WrAddr_cole, Q => 
        \SD_WrAddr_col[8]_net_1\);
    
    \temp_w[1]\ : DFN1C0
      port map(D => \temp_w_n1_0_i_0\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \temp_w[1]_net_1\);
    
    \SD_wrAddr_row_RNO[12]\ : XA1
      port map(A => N237_0, B => ADD_13x13_medium_area_I49_Y_0_0, 
        C => un7_sdram_enreg, Y => \SD_wrAddr_row_6[12]\);
    
    \addr_RNO_0[1]\ : OA1A
      port map(A => \SD_wrAddr_row[1]_net_1\, B => N_191, C => 
        N_303, Y => \addr_11_0_0_0[1]\);
    
    WFifo_re_RNO_0 : OR3A
      port map(A => \Z\\SDRAM_wr_0_wr_state_[2]\\\, B => 
        \Z\\SDRAM_wr_0_wr_state_[0]\\\, C => un1_cs_n7_4_i_0_a7_0, 
        Y => un1_cs_n7_4_i_0_a7_1);
    
    \addr_RNO[1]\ : OR3C
      port map(A => \addr_11_0_0_0[1]\, B => N_304, C => N_249_i, 
        Y => \addr_11[1]\);
    
    \SD_rdAddr_col[7]\ : DFN1E1C0
      port map(D => N_542, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => SD_rdAddr_cole, Q => 
        \SD_rdAddr_col[7]_net_1\);
    
    ras_n : DFN1P0
      port map(D => ras_n_5, CLK => PLL_Test1_0_Sys_66M_Clk, PRE
         => PLL_Test1_0_SysRst_O, Q => SD_ras_n_c);
    
    \addr[3]\ : DFN1C0
      port map(D => N_164_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \SD_addr_c[3]\);
    
    \SD_rdAddr_col[4]\ : DFN1E1C0
      port map(D => N_540, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => SD_rdAddr_cole, Q => 
        \SD_rdAddr_col[4]_net_1\);
    
    \addr_RNO[11]\ : NOR3
      port map(A => N_340, B => N_342, C => N_633, Y => N_176);
    
    un1_SD_wrAddr_row_ADD_13x13_medium_area_I10_Y : NOR2B
      port map(A => N153, B => \SD_wrAddr_row[1]_net_1\, Y => 
        N215_0);
    
    \addr_RNO_4[6]\ : OR3A
      port map(A => N_186, B => N_371, C => 
        \SD_rdAddr_col[6]_net_1\, Y => \addr_RNO_4[6]_net_1\);
    
    cas_n_RNO : OAI1
      port map(A => N_353_2, B => cas_n_4_6_0_a7_1_0, C => 
        cas_n_4_6_0_0_1, Y => cas_n_4);
    
    \addr_RNO_0[3]\ : NOR3C
      port map(A => \addr_RNO_2[3]_net_1\, B => 
        \addr_RNO_3[3]_net_1\, C => \addr_11_0_i_0[3]\, Y => 
        \addr_11_0_i_2[3]\);
    
    un1_SD_rdAddr_row_ADD_13x13_medium_area_I14_Y_0 : OR2B
      port map(A => \SD_rdAddr_row[3]_net_1\, B => 
        \SD_rdAddr_row[2]_net_1\, Y => 
        ADD_13x13_medium_area_I14_Y_0_0);
    
    \SD_WrAddr_col_RNI2S3F[6]\ : NOR2A
      port map(A => \SD_WrAddr_col[6]_net_1\, B => N_196, Y => 
        N_199);
    
    temp_w_n2_0_i_0 : XA1
      port map(A => N_207, B => \temp_w[2]_net_1\, C => N_191, Y
         => \temp_w_n2_0_i_0\);
    
    \SD_WrAddr_col_RNO[5]\ : NOR3B
      port map(A => N_196, B => N_255, C => un1_sdram_enreg_2, Y
         => N_11_i_0);
    
    rdrow_end_RNO_2 : NOR3
      port map(A => \SD_rdAddr_col[5]_net_1\, B => 
        \SD_rdAddr_col[4]_net_1\, C => \SD_rdAddr_col[10]_net_1\, 
        Y => un4lt10_i_a2_0_a7_3);
    
    \SD_wrAddr_row_RNI0TRI[1]\ : NOR3A
      port map(A => sd_wraddr_row20_0_a7_2, B => 
        \SD_wrAddr_row[3]_net_1\, C => \SD_wrAddr_row[1]_net_1\, 
        Y => sd_wraddr_row20_0_a7_7);
    
    \addr_RNO[2]\ : NOR3C
      port map(A => \addr_11_0_i_0[2]\, B => N_372, C => 
        \addr_11_0_i_2[2]\, Y => N_162_i_0);
    
    \SD_rdAddr_row[1]\ : DFN1C0
      port map(D => \SD_rdAddr_row_6[1]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \SD_rdAddr_row[1]_net_1\);
    
    \SD_rdAddr_col_RNO_0[7]\ : AOI1
      port map(A => \SD_rdAddr_col[6]_net_1\, B => N_197, C => 
        \SD_rdAddr_col[7]_net_1\, Y => N_297);
    
    \SD_rdAddr_row[6]\ : DFN1C0
      port map(D => \SD_rdAddr_row_6[6]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \SD_rdAddr_row[6]_net_1\);
    
    \addr_RNO_0[9]\ : NOR3C
      port map(A => \addr_RNO_2[9]_net_1\, B => N_253, C => 
        \addr_RNO_4[9]_net_1\, Y => \addr_11_i_0_2[9]\);
    
    un1_SD_rdAddr_row_ADD_13x13_medium_area_I22_Y : AO1B
      port map(A => ADD_13x13_medium_area_I22_un1_Y_1_0, B => 
        N245, C => sd_rdaddr_row18_i, Y => N237);
    
    \SD_rdAddr_col[5]\ : DFN1E1C0
      port map(D => N_35, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => SD_rdAddr_cole, Q => 
        \SD_rdAddr_col[5]_net_1\);
    
    \addr_RNO_1[3]\ : OR3A
      port map(A => N_186, B => N_371, C => 
        \SD_rdAddr_col[3]_net_1\, Y => \addr_RNO_1[3]_net_1\);
    
    \addr_11_i_0_a2_1[9]\ : OR2B
      port map(A => N_198, B => \Z\\Sdram_ini_0_ini_state_[2]\\\, 
        Y => N_384);
    
    \SD_WrAddr_col_RNID9611_0[10]\ : NOR2A
      port map(A => \un1_sd_wraddr_row8_i_0[12]\, B => N_239, Y
         => \un1_sd_wraddr_row8_i_1[12]\);
    
    \SD_wrAddr_row[4]\ : DFN1C0
      port map(D => \SD_wrAddr_row_6[4]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \SD_wrAddr_row[4]_net_1\);
    
    \SD_rdAddr_col[9]\ : DFN1E1C0
      port map(D => N_544, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => SD_rdAddr_cole, Q => 
        \SD_rdAddr_col[9]_net_1\);
    
    \dqm_1_RNO_0[0]\ : NOR3A
      port map(A => \Z\\SDram_rd_0_rd_state_[2]\\\, B => 
        \Z\\SDram_rd_0_rd_state_[1]\\\, C => N_221, Y => N_263);
    
    \addr_RNO_0[11]\ : AOI1
      port map(A => N_384, B => \SD_addr_c[11]\, C => N_343_1, Y
         => N_340);
    
    \addr_RNO_9[10]\ : NOR2A
      port map(A => \SD_wrAddr_row[10]_net_1\, B => 
        \Z\\SDRAM_wr_0_wr_state_[2]\\\, Y => N_225);
    
    \SD_rdAddr_col[10]\ : DFN1C0
      port map(D => \SD_rdAddr_col_RNO[10]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \SD_rdAddr_col[10]_net_1\);
    
    un1_SD_rdAddr_row_ADD_13x13_medium_area_I15_Y_1 : NOR3C
      port map(A => \SD_rdAddr_row[6]_net_1\, B => 
        \SD_rdAddr_row[7]_net_1\, C => N253_0, Y => 
        ADD_13x13_medium_area_I15_Y_1_0);
    
    ras_n_5_7_0_o4_0 : OR2A
      port map(A => \Z\\SDram_rd_0_rd_state_[1]\\\, B => 
        \Z\\SDram_rd_0_rd_state_[0]\\\, Y => N_190);
    
    un1_SD_wrAddr_row_ADD_13x13_medium_area_I32_Y : NOR2B
      port map(A => N256_0, B => N253, Y => N258_0);
    
    wrrow_end : DFN1E1C0
      port map(D => \SD_WrAddr_col[9]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => N_4, Q => Sdram_cmd_0_wrrow_end);
    
    \SD_wrAddr_row_RNO[3]\ : XA1A
      port map(A => \SD_wrAddr_row[3]_net_1\, B => I37_un1_Y_0, C
         => un7_sdram_enreg, Y => \SD_wrAddr_row_6[3]\);
    
    \SD_wrAddr_row_RNO[5]\ : XA1A
      port map(A => \SD_wrAddr_row[5]_net_1\, B => I36_un1_Y_0, C
         => un7_sdram_enreg, Y => \SD_wrAddr_row_6[5]\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3;
use proasic3.all;

entity Sdram_ini is

    port( \Z\\Sdram_ini_0_ini_state_[2]\\\ : out   std_logic;
          \Z\\Sdram_ini_0_ini_state_[1]\\\ : out   std_logic;
          \Z\\Sdram_ini_0_ini_state_[0]\\\ : out   std_logic;
          PLL_Test1_0_SysRst_O             : in    std_logic;
          PLL_Test1_0_Sys_66M_Clk          : in    std_logic;
          Sdram_ctl_v2_0_SD_iniEn          : in    std_logic;
          Sdram_ini_0_Sd_iniOK             : out   std_logic;
          Sdram_ini_0_Sd_iniOK_i           : out   std_logic
        );

end Sdram_ini;

architecture DEF_ARCH of Sdram_ini is 

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component INV
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OAI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XNOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XAI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component AO1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NOR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \pr_state_ns_0_a3_4_a2_1[0]\, \pr_state[0]_net_1\, 
        \pr_state[1]_net_1\, \pr_state_RNI0ICC[2]_net_1\, 
        \pr_state_ns_0_i_0[5]\, trc_nume, pr_state_tr10_i_a2_0, 
        \counter_200[12]_net_1\, \counter_200[13]_net_1\, 
        \pr_state_ns_0_0_a2_0_0[1]\, N_195_1, N_49, 
        pr_state_tr7_i_a2_0, \trc_num[0]_net_1\, 
        \trc_num[1]_net_1\, \pr_state_ns_0_0_a2_1_0[1]\, 
        \refresh_timer[3]_net_1\, \refresh_timer_i[2]\, 
        pr_state_tr10_i_a2_0_1, \counter_200[7]_net_1\, 
        \counter_200[8]_net_1\, pr_state_tr10_i_a2_0_0, 
        \counter_200[5]_net_1\, \counter_200[6]_net_1\, N_12_i_0, 
        \counter_200[0]_net_1\, \counter_200[1]_net_1\, 
        \pr_state[5]_net_1\, N_14_i_0, N_47, 
        \counter_200[2]_net_1\, N_17, N_48, 
        \counter_200[3]_net_1\, \counter_200_RNO[4]_net_1\, N_110, 
        N_51, \counter_200_RNO[5]_net_1\, 
        \counter_200_RNO[6]_net_1\, N_52, N_26, N_53, 
        \counter_200_RNO[8]_net_1\, N_54, 
        \ini_state_RNO[0]_net_1\, \pr_state[3]_net_1\, N_9, N_144, 
        \pr_state_ns[2]\, N_41, \refresh_timer[0]_net_1\, 
        \refresh_timer[1]_net_1\, N_8, N_20, N_40, trc_num_n3, 
        N_21, \trc_num[2]_net_1\, \trc_num[3]_net_1\, 
        \pr_state_RNO[2]_net_1\, counter_200_n0, 
        \counter_200[4]_net_1\, counter_200_n9, 
        \counter_200[9]_net_1\, N_56, counter_200_n10, 
        \counter_200[10]_net_1\, N_95, counter_200_n11, 
        \counter_200[11]_net_1\, N_94, counter_200_n12, N_59, 
        counter_200_n13, N_92, counter_200_n14, 
        \counter_200[14]_net_1\, N_193, \pr_state_ns[0]\, N_91, 
        N_57, N_87, N_89, \pr_state_RNO[1]_net_1\, 
        \pr_state_ns[1]\, N_194, \pr_state[2]_net_1\, 
        refresh_timer_n0, N_25_i, N_24_i, N_22, N_10, 
        \ini_state_RNO[2]_net_1\, N_27_i_i_0, N_35, 
        \Sdram_ini_0_Sd_iniOK\, \GND\, \VCC\, GND_0, VCC_0
         : std_logic;

begin 

    Sdram_ini_0_Sd_iniOK <= \Sdram_ini_0_Sd_iniOK\;

    \trc_num_RNO[0]\ : XOR2
      port map(A => trc_nume, B => \trc_num[0]_net_1\, Y => 
        N_25_i);
    
    \counter_200_RNO[14]\ : XA1A
      port map(A => \counter_200[14]_net_1\, B => N_193, C => 
        \pr_state[5]_net_1\, Y => counter_200_n14);
    
    \counter_200_RNO[9]\ : XA1A
      port map(A => \counter_200[9]_net_1\, B => N_56, C => 
        \pr_state[5]_net_1\, Y => counter_200_n9);
    
    \counter_200_RNO[11]\ : XA1A
      port map(A => \counter_200[11]_net_1\, B => N_94, C => 
        \pr_state[5]_net_1\, Y => counter_200_n11);
    
    \refresh_timer_RNIUVOE[1]\ : NOR3
      port map(A => \refresh_timer[0]_net_1\, B => 
        \refresh_timer[1]_net_1\, C => 
        \pr_state_ns_0_0_a2_1_0[1]\, Y => N_144);
    
    \pr_state_RNI0ICC[2]\ : OR2
      port map(A => trc_nume, B => \pr_state[2]_net_1\, Y => 
        \pr_state_RNI0ICC[2]_net_1\);
    
    \counter_200[2]\ : DFN1C0
      port map(D => N_14_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \counter_200[2]_net_1\);
    
    \counter_200_RNIU3EN1[12]\ : OA1B
      port map(A => N_87, B => pr_state_tr10_i_a2_0, C => N_89, Y
         => N_91);
    
    \counter_200_RNO[1]\ : XA1
      port map(A => \counter_200[0]_net_1\, B => 
        \counter_200[1]_net_1\, C => \pr_state[5]_net_1\, Y => 
        N_12_i_0);
    
    \pr_state_RNO_0[5]\ : OR3
      port map(A => \pr_state[0]_net_1\, B => \pr_state[1]_net_1\, 
        C => \pr_state_RNI0ICC[2]_net_1\, Y => 
        \pr_state_ns_0_a3_4_a2_1[0]\);
    
    \pr_state_RNO_0[4]\ : NOR2A
      port map(A => N_195_1, B => N_49, Y => 
        \pr_state_ns_0_0_a2_0_0[1]\);
    
    \trc_num_RNIN5D8[3]\ : OR2A
      port map(A => \trc_num[3]_net_1\, B => \trc_num[2]_net_1\, 
        Y => N_40);
    
    \refresh_timer[0]\ : DFN1C0
      port map(D => refresh_timer_n0, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \refresh_timer[0]_net_1\);
    
    \counter_200_RNIQTHG[4]\ : NOR3B
      port map(A => \counter_200[3]_net_1\, B => 
        \counter_200[4]_net_1\, C => N_48, Y => N_51);
    
    \pr_state_RNO_1[4]\ : OR2B
      port map(A => \pr_state[2]_net_1\, B => 
        Sdram_ctl_v2_0_SD_iniEn, Y => N_194);
    
    \counter_200_RNI5P6N[6]\ : NOR2B
      port map(A => \counter_200[6]_net_1\, B => N_52, Y => N_53);
    
    \counter_200_RNIJIT9[2]\ : OR2A
      port map(A => \counter_200[2]_net_1\, B => N_47, Y => N_48);
    
    \refresh_timer_RNO_0[3]\ : NOR2
      port map(A => \refresh_timer_i[2]\, B => N_20, Y => N_22);
    
    \refresh_timer[3]\ : DFN1C0
      port map(D => N_10, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \refresh_timer[3]_net_1\);
    
    \counter_200_RNO[3]\ : XA1A
      port map(A => N_48, B => \counter_200[3]_net_1\, C => 
        \pr_state[5]_net_1\, Y => N_17);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \ini_state_RNO[2]\ : OR2
      port map(A => \pr_state[3]_net_1\, B => \pr_state[0]_net_1\, 
        Y => \ini_state_RNO[2]_net_1\);
    
    \counter_200_RNIQ5MT[5]\ : OA1B
      port map(A => pr_state_tr10_i_a2_0_0, B => 
        pr_state_tr10_i_a2_0_1, C => N_57, Y => N_87);
    
    \trc_num_RNIARPG[1]\ : NOR2
      port map(A => pr_state_tr7_i_a2_0, B => N_40, Y => N_49);
    
    \counter_200_RNIK4ST[8]\ : OR2B
      port map(A => \counter_200[8]_net_1\, B => N_54, Y => N_56);
    
    \counter_200[4]\ : DFN1C0
      port map(D => \counter_200_RNO[4]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \counter_200[4]_net_1\);
    
    \refresh_timer[2]\ : DFN1P0
      port map(D => N_8, CLK => PLL_Test1_0_Sys_66M_Clk, PRE => 
        PLL_Test1_0_SysRst_O, Q => \refresh_timer_i[2]\);
    
    Sd_iniOK_RNI7HH2 : INV
      port map(A => \Sdram_ini_0_Sd_iniOK\, Y => 
        Sdram_ini_0_Sd_iniOK_i);
    
    \trc_num_RNIJLC8_0[1]\ : OR2
      port map(A => \trc_num[0]_net_1\, B => \trc_num[1]_net_1\, 
        Y => pr_state_tr7_i_a2_0);
    
    \counter_200_RNO[0]\ : NOR2A
      port map(A => \pr_state[5]_net_1\, B => 
        \counter_200[0]_net_1\, Y => counter_200_n0);
    
    \trc_num[0]\ : DFN1C0
      port map(D => N_25_i, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \trc_num[0]_net_1\);
    
    \refresh_timer[1]\ : DFN1C0
      port map(D => N_41, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \refresh_timer[1]_net_1\);
    
    \counter_200_RNO_0[11]\ : OR3B
      port map(A => \counter_200[9]_net_1\, B => 
        \counter_200[10]_net_1\, C => N_56, Y => N_94);
    
    \counter_200[14]\ : DFN1C0
      port map(D => counter_200_n14, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \counter_200[14]_net_1\);
    
    \counter_200[13]\ : DFN1C0
      port map(D => counter_200_n13, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \counter_200[13]_net_1\);
    
    \pr_state_RNO[5]\ : OAI1
      port map(A => N_91, B => \pr_state_ns_0_a3_4_a2_1[0]\, C
         => Sdram_ctl_v2_0_SD_iniEn, Y => \pr_state_ns[0]\);
    
    \pr_state[3]\ : DFN1C0
      port map(D => \pr_state_ns[2]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \pr_state[3]_net_1\);
    
    \ini_state[1]\ : DFN1C0
      port map(D => \pr_state_RNI0ICC[2]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \Z\\Sdram_ini_0_ini_state_[1]\\\);
    
    \refresh_timer_RNIT7C7[1]\ : OR2B
      port map(A => \refresh_timer[1]_net_1\, B => 
        \refresh_timer[0]_net_1\, Y => N_20);
    
    \refresh_timer_RNI1OC7[3]\ : OR2
      port map(A => \refresh_timer[3]_net_1\, B => 
        \refresh_timer_i[2]\, Y => \pr_state_ns_0_0_a2_1_0[1]\);
    
    \pr_state_RNO_0[0]\ : OA1
      port map(A => \pr_state[0]_net_1\, B => trc_nume, C => 
        Sdram_ctl_v2_0_SD_iniEn, Y => \pr_state_ns_0_i_0[5]\);
    
    \counter_200_RNIB31D[12]\ : OR2
      port map(A => \counter_200[12]_net_1\, B => 
        \counter_200[13]_net_1\, Y => pr_state_tr10_i_a2_0);
    
    \refresh_timer_RNO[3]\ : XA1
      port map(A => N_22, B => \refresh_timer[3]_net_1\, C => 
        \pr_state[0]_net_1\, Y => N_10);
    
    \pr_state[2]\ : DFN1C0
      port map(D => \pr_state_RNO[2]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \pr_state[2]_net_1\);
    
    \pr_state_RNO[0]\ : OA1A
      port map(A => N_144, B => trc_nume, C => 
        \pr_state_ns_0_i_0[5]\, Y => N_9);
    
    \counter_200_RNO[13]\ : XA1A
      port map(A => \counter_200[13]_net_1\, B => N_92, C => 
        \pr_state[5]_net_1\, Y => counter_200_n13);
    
    \counter_200_RNIBRK6[5]\ : OR2
      port map(A => \counter_200[5]_net_1\, B => 
        \counter_200[6]_net_1\, Y => pr_state_tr10_i_a2_0_0);
    
    \counter_200_RNIF9SJ[5]\ : NOR2B
      port map(A => \counter_200[5]_net_1\, B => N_51, Y => N_52);
    
    \trc_num_RNO[2]\ : XNOR2
      port map(A => \trc_num[2]_net_1\, B => N_21, Y => 
        N_27_i_i_0);
    
    \refresh_timer_RNO[2]\ : XAI1
      port map(A => N_20, B => \refresh_timer_i[2]\, C => 
        \pr_state[0]_net_1\, Y => N_8);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \counter_200_RNO_0[10]\ : OR2A
      port map(A => \counter_200[9]_net_1\, B => N_56, Y => N_95);
    
    \trc_num_RNIJLC8[1]\ : OR2B
      port map(A => \trc_num[1]_net_1\, B => \trc_num[0]_net_1\, 
        Y => N_21);
    
    \counter_200[8]\ : DFN1C0
      port map(D => \counter_200_RNO[8]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \counter_200[8]_net_1\);
    
    \pr_state_RNO[4]\ : AO1B
      port map(A => \pr_state_ns_0_0_a2_0_0[1]\, B => N_144, C
         => N_194, Y => \pr_state_ns[1]\);
    
    \pr_state_RNO[1]\ : NOR2B
      port map(A => N_91, B => Sdram_ctl_v2_0_SD_iniEn, Y => 
        \pr_state_RNO[1]_net_1\);
    
    \counter_200_RNO[5]\ : XA1
      port map(A => N_51, B => \counter_200[5]_net_1\, C => 
        \pr_state[5]_net_1\, Y => \counter_200_RNO[5]_net_1\);
    
    \counter_200[11]\ : DFN1C0
      port map(D => counter_200_n11, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \counter_200[11]_net_1\);
    
    \counter_200[12]\ : DFN1C0
      port map(D => counter_200_n12, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \counter_200[12]_net_1\);
    
    \pr_state[0]\ : DFN1C0
      port map(D => N_9, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \pr_state[0]_net_1\);
    
    \counter_200_RNI9LOK1[12]\ : OR2B
      port map(A => \counter_200[12]_net_1\, B => N_59, Y => N_92);
    
    \counter_200[10]\ : DFN1C0
      port map(D => counter_200_n10, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \counter_200[10]_net_1\);
    
    \counter_200[0]\ : DFN1C0
      port map(D => counter_200_n0, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \counter_200[0]_net_1\);
    
    \pr_state_RNO[2]\ : NOR2B
      port map(A => \pr_state[1]_net_1\, B => 
        Sdram_ctl_v2_0_SD_iniEn, Y => \pr_state_RNO[2]_net_1\);
    
    \counter_200_RNO[10]\ : XA1A
      port map(A => \counter_200[10]_net_1\, B => N_95, C => 
        \pr_state[5]_net_1\, Y => counter_200_n10);
    
    \trc_num[1]\ : DFN1E1C0
      port map(D => N_24_i, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => trc_nume, Q => 
        \trc_num[1]_net_1\);
    
    \counter_200[9]\ : DFN1C0
      port map(D => counter_200_n9, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \counter_200[9]_net_1\);
    
    \ini_state_RNO[0]\ : OR3
      port map(A => \pr_state[3]_net_1\, B => \pr_state[1]_net_1\, 
        C => trc_nume, Y => \ini_state_RNO[0]_net_1\);
    
    \trc_num[2]\ : DFN1E1C0
      port map(D => N_27_i_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => trc_nume, Q => 
        \trc_num[2]_net_1\);
    
    \ini_state[2]\ : DFN1C0
      port map(D => \ini_state_RNO[2]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \Z\\Sdram_ini_0_ini_state_[2]\\\);
    
    \counter_200[6]\ : DFN1C0
      port map(D => \counter_200_RNO[6]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \counter_200[6]_net_1\);
    
    \pr_state[4]\ : DFN1C0
      port map(D => \pr_state_ns[1]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => trc_nume);
    
    \ini_state[0]\ : DFN1C0
      port map(D => \ini_state_RNO[0]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \Z\\Sdram_ini_0_ini_state_[0]\\\);
    
    \counter_200_RNO_0[14]\ : OR2A
      port map(A => \counter_200[13]_net_1\, B => N_92, Y => 
        N_193);
    
    Sd_iniOK : DFN1C0
      port map(D => N_35, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Sdram_ini_0_Sd_iniOK\);
    
    \counter_200_RNO[4]\ : NOR3A
      port map(A => \pr_state[5]_net_1\, B => N_110, C => N_51, Y
         => \counter_200_RNO[4]_net_1\);
    
    \counter_200_RNIK38E1[11]\ : NOR2
      port map(A => N_57, B => N_56, Y => N_59);
    
    \counter_200_RNO_0[4]\ : OA1C
      port map(A => \counter_200[3]_net_1\, B => N_48, C => 
        \counter_200[4]_net_1\, Y => N_110);
    
    \counter_200[3]\ : DFN1C0
      port map(D => N_17, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \counter_200[3]_net_1\);
    
    \trc_num[3]\ : DFN1E1C0
      port map(D => trc_num_n3, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => trc_nume, Q => 
        \trc_num[3]_net_1\);
    
    \pr_state_RNIJ2SD[0]\ : NOR2B
      port map(A => \pr_state[0]_net_1\, B => 
        Sdram_ctl_v2_0_SD_iniEn, Y => N_195_1);
    
    \counter_200_RNO[6]\ : XA1
      port map(A => N_52, B => \counter_200[6]_net_1\, C => 
        \pr_state[5]_net_1\, Y => \counter_200_RNO[6]_net_1\);
    
    \counter_200_RNO[8]\ : XA1
      port map(A => N_54, B => \counter_200[8]_net_1\, C => 
        \pr_state[5]_net_1\, Y => \counter_200_RNO[8]_net_1\);
    
    \counter_200_RNIFBL6[7]\ : OR2
      port map(A => \counter_200[7]_net_1\, B => 
        \counter_200[8]_net_1\, Y => pr_state_tr10_i_a2_0_1);
    
    \pr_state[1]\ : DFN1C0
      port map(D => \pr_state_RNO[1]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \pr_state[1]_net_1\);
    
    Sd_iniOK_RNO : OR2
      port map(A => \Sdram_ini_0_Sd_iniOK\, B => 
        \pr_state[3]_net_1\, Y => N_35);
    
    \counter_200_RNO[12]\ : XA1
      port map(A => \counter_200[12]_net_1\, B => N_59, C => 
        \pr_state[5]_net_1\, Y => counter_200_n12);
    
    \counter_200_RNO[7]\ : XA1
      port map(A => N_53, B => \counter_200[7]_net_1\, C => 
        \pr_state[5]_net_1\, Y => N_26);
    
    \counter_200_RNI0VBG[11]\ : OR3C
      port map(A => \counter_200[9]_net_1\, B => 
        \counter_200[10]_net_1\, C => \counter_200[11]_net_1\, Y
         => N_57);
    
    \counter_200[1]\ : DFN1C0
      port map(D => N_12_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \counter_200[1]_net_1\);
    
    \pr_state[5]\ : DFN1P0
      port map(D => \pr_state_ns[0]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, PRE => PLL_Test1_0_SysRst_O, Q
         => \pr_state[5]_net_1\);
    
    \counter_200_RNI1JJ6[1]\ : OR2B
      port map(A => \counter_200[1]_net_1\, B => 
        \counter_200[0]_net_1\, Y => N_47);
    
    \refresh_timer_RNO[1]\ : XA1
      port map(A => \refresh_timer[0]_net_1\, B => 
        \refresh_timer[1]_net_1\, C => \pr_state[0]_net_1\, Y => 
        N_41);
    
    \counter_200[7]\ : DFN1C0
      port map(D => N_26, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \counter_200[7]_net_1\);
    
    \trc_num_RNO[1]\ : XOR2
      port map(A => \trc_num[1]_net_1\, B => \trc_num[0]_net_1\, 
        Y => N_24_i);
    
    \pr_state_RNO[3]\ : NOR3C
      port map(A => N_49, B => N_195_1, C => N_144, Y => 
        \pr_state_ns[2]\);
    
    \counter_200_RNISCHQ[7]\ : NOR2B
      port map(A => \counter_200[7]_net_1\, B => N_53, Y => N_54);
    
    \refresh_timer_RNO[0]\ : NOR2A
      port map(A => \pr_state[0]_net_1\, B => 
        \refresh_timer[0]_net_1\, Y => refresh_timer_n0);
    
    \counter_200_RNIPQMC[14]\ : OR2B
      port map(A => \pr_state[5]_net_1\, B => 
        \counter_200[14]_net_1\, Y => N_89);
    
    \counter_200[5]\ : DFN1C0
      port map(D => \counter_200_RNO[5]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \counter_200[5]_net_1\);
    
    \counter_200_RNO[2]\ : XA1A
      port map(A => N_47, B => \counter_200[2]_net_1\, C => 
        \pr_state[5]_net_1\, Y => N_14_i_0);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    \trc_num_RNO[3]\ : AX1
      port map(A => N_21, B => \trc_num[2]_net_1\, C => 
        \trc_num[3]_net_1\, Y => trc_num_n3);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3;
use proasic3.all;

entity SDram_rd is

    port( \Z\\SDram_rd_0_rd_state_[2]\\\ : out   std_logic;
          \Z\\SDram_rd_0_rd_state_[1]\\\ : out   std_logic;
          \Z\\SDram_rd_0_rd_state_[0]\\\ : out   std_logic;
          Sdram_ctl_v2_0_SD_rdEn_i       : in    std_logic;
          PLL_Test1_0_SysRst_O           : in    std_logic;
          PLL_Test1_0_Sys_66M_Clk        : in    std_logic;
          SDram_rd_0_SD_RdOK             : out   std_logic;
          Sdram_ctl_v2_0_SD_rdEn         : in    std_logic;
          Sdram_cmd_0_rdrow_end          : in    std_logic;
          Sdram_ctl_v2_0_SD_rdEN_noact   : in    std_logic
        );

end SDram_rd;

architecture DEF_ARCH of SDram_rd is 

  component OR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component XNOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \pr_state_ns_0_a2_0_0[1]\, 
        \rd_state_9_0_i_a2_0_a2_0[2]\, \pr_state[1]_net_1\, 
        \pr_state[0]_net_1\, \rd_state_9_0_i_a2_0_a2_0[1]\, 
        \pr_state[4]_net_1\, \pr_state[6]_net_1\, N_22, 
        \pr_state[3]_net_1\, \temp_i[1]\, N_26_i_i_0, 
        \rd_state_RNO[1]_net_1\, \rd_state_RNO[2]_net_1\, 
        \pr_state[5]_net_1\, \rd_state_RNO[0]_net_1\, N_51, 
        \pr_state_ns[5]\, N_49, rd_ok_0_sqmuxa, \temp[2]_net_1\, 
        N_76_i, N_43, \pr_state[2]_net_1\, 
        \pr_state_RNO[5]_net_1\, \pr_state_RNO_0[3]\, N_18, 
        \temp[0]_net_1\, N_24, N_20, \pr_state_ns[1]\, N_101, 
        \pr_state[7]_net_1\, N_42, \GND\, \VCC\, GND_0, VCC_0
         : std_logic;

begin 


    \rd_state_RNO[2]\ : OR3
      port map(A => \pr_state[3]_net_1\, B => \pr_state[5]_net_1\, 
        C => \rd_state_9_0_i_a2_0_a2_0[2]\, Y => 
        \rd_state_RNO[2]_net_1\);
    
    rd_ok_RNO : NOR3C
      port map(A => \temp[2]_net_1\, B => \temp_i[1]\, C => 
        \pr_state[3]_net_1\, Y => rd_ok_0_sqmuxa);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \rd_state_RNO[0]\ : OR3
      port map(A => \pr_state[0]_net_1\, B => N_51, C => 
        \pr_state[3]_net_1\, Y => \rd_state_RNO[0]_net_1\);
    
    temp_n0_0_i : NOR2
      port map(A => \temp[0]_net_1\, B => N_24, Y => N_18);
    
    \pr_state_RNO[6]\ : AO1B
      port map(A => \pr_state_ns_0_a2_0_0[1]\, B => N_49, C => 
        N_101, Y => \pr_state_ns[1]\);
    
    \rd_state[2]\ : DFN1C0
      port map(D => \rd_state_RNO[2]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \Z\\SDram_rd_0_rd_state_[2]\\\);
    
    \pr_state_RNO_0[6]\ : NOR2
      port map(A => Sdram_ctl_v2_0_SD_rdEN_noact, B => 
        Sdram_cmd_0_rdrow_end, Y => \pr_state_ns_0_a2_0_0[1]\);
    
    \pr_state_RNO[5]\ : NOR2B
      port map(A => Sdram_ctl_v2_0_SD_rdEn, B => N_51, Y => 
        \pr_state_RNO[5]_net_1\);
    
    \pr_state[3]\ : DFN1C0
      port map(D => \pr_state_RNO_0[3]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \pr_state[3]_net_1\);
    
    \temp[1]\ : DFN1P0
      port map(D => N_20, CLK => PLL_Test1_0_Sys_66M_Clk, PRE => 
        PLL_Test1_0_SysRst_O, Q => \temp_i[1]\);
    
    \pr_state_RNO_1[6]\ : OR2B
      port map(A => Sdram_ctl_v2_0_SD_rdEn, B => 
        \pr_state[0]_net_1\, Y => N_101);
    
    \pr_state[2]\ : DFN1C0
      port map(D => \pr_state_ns[5]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \pr_state[2]_net_1\);
    
    \pr_state_RNO[0]\ : NOR2B
      port map(A => Sdram_ctl_v2_0_SD_rdEn, B => 
        \pr_state[1]_net_1\, Y => N_43);
    
    \temp[2]\ : DFN1C0
      port map(D => N_22, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \temp[2]_net_1\);
    
    \pr_state[7]\ : DFN1P0
      port map(D => Sdram_ctl_v2_0_SD_rdEn_i, CLK => 
        PLL_Test1_0_Sys_66M_Clk, PRE => PLL_Test1_0_SysRst_O, Q
         => \pr_state[7]_net_1\);
    
    \rd_state[0]\ : DFN1C0
      port map(D => \rd_state_RNO[0]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \Z\\SDram_rd_0_rd_state_[0]\\\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \pr_state_RNO[4]\ : NOR2B
      port map(A => Sdram_ctl_v2_0_SD_rdEn, B => 
        \pr_state[6]_net_1\, Y => N_76_i);
    
    \pr_state_RNO[1]\ : NOR2B
      port map(A => Sdram_cmd_0_rdrow_end, B => N_49, Y => N_42);
    
    \pr_state[0]\ : DFN1C0
      port map(D => N_43, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \pr_state[0]_net_1\);
    
    temp_n2_0_i_x2 : XNOR2
      port map(A => \temp[2]_net_1\, B => \temp[0]_net_1\, Y => 
        N_26_i_i_0);
    
    \pr_state_RNO[2]\ : NOR3B
      port map(A => Sdram_ctl_v2_0_SD_rdEN_noact, B => N_49, C
         => Sdram_cmd_0_rdrow_end, Y => \pr_state_ns[5]\);
    
    rd_ok : DFN1C0
      port map(D => rd_ok_0_sqmuxa, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => SDram_rd_0_SD_RdOK);
    
    \temp[0]\ : DFN1C0
      port map(D => N_18, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \temp[0]_net_1\);
    
    \pr_state_RNIG4M6[7]\ : NOR2B
      port map(A => Sdram_ctl_v2_0_SD_rdEn, B => 
        \pr_state[7]_net_1\, Y => N_49);
    
    \pr_state_RNIKG76[2]\ : OR2
      port map(A => \pr_state[4]_net_1\, B => \pr_state[2]_net_1\, 
        Y => N_51);
    
    \rd_state[1]\ : DFN1C0
      port map(D => \rd_state_RNO[1]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \Z\\SDram_rd_0_rd_state_[1]\\\);
    
    \pr_state[4]\ : DFN1C0
      port map(D => N_76_i, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \pr_state[4]_net_1\);
    
    \pr_state[6]\ : DFN1C0
      port map(D => \pr_state_ns[1]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \pr_state[6]_net_1\);
    
    \rd_state_RNO_0[1]\ : OR2
      port map(A => \pr_state[4]_net_1\, B => \pr_state[6]_net_1\, 
        Y => \rd_state_9_0_i_a2_0_a2_0[1]\);
    
    \pr_state[1]\ : DFN1C0
      port map(D => N_42, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \pr_state[1]_net_1\);
    
    \pr_state[5]\ : DFN1C0
      port map(D => \pr_state_RNO[5]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \pr_state[5]_net_1\);
    
    temp_n1_0_i : XO1
      port map(A => \temp[0]_net_1\, B => \temp_i[1]\, C => N_24, 
        Y => N_20);
    
    temp_n0_0_i_o2 : AO1B
      port map(A => \temp_i[1]\, B => \temp[2]_net_1\, C => 
        \pr_state[3]_net_1\, Y => N_24);
    
    \rd_state_RNO_0[2]\ : OR2
      port map(A => \pr_state[1]_net_1\, B => \pr_state[0]_net_1\, 
        Y => \rd_state_9_0_i_a2_0_a2_0[2]\);
    
    \pr_state_RNO[3]\ : OA1
      port map(A => \pr_state[3]_net_1\, B => \pr_state[5]_net_1\, 
        C => Sdram_ctl_v2_0_SD_rdEn, Y => \pr_state_RNO_0[3]\);
    
    temp_n2_0_i : NOR3A
      port map(A => \pr_state[3]_net_1\, B => \temp_i[1]\, C => 
        N_26_i_i_0, Y => N_22);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    \rd_state_RNO[1]\ : OR3
      port map(A => \rd_state_9_0_i_a2_0_a2_0[1]\, B => 
        \pr_state[1]_net_1\, C => \pr_state[0]_net_1\, Y => 
        \rd_state_RNO[1]_net_1\);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3;
use proasic3.all;

entity WaveGenSingleZ11 is

    port( CMOS_DrvX_0_LVDSen_2    : in    std_logic;
          CMOS_DrvX_0_LVDSen_1    : in    std_logic;
          lvdsFifoRowRdOut        : out   std_logic;
          lvdsFifoRowRdOut_i      : out   std_logic;
          PLL_Test1_0_SysRst_O    : in    std_logic;
          PLL_Test1_0_Sys_66M_Clk : in    std_logic
        );

end WaveGenSingleZ11;

architecture DEF_ARCH of WaveGenSingleZ11 is 

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NOR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OAI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component INV
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1E
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component XA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component XA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component AOI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \PrState_0[1]_net_1\, N_8, \PrState_ns_0_i_0_a3_0[2]\, 
        N_242, \PrState[2]_net_1\, N_166, 
        \PrState_ns_0_i_0_a3_0_0[2]\, \CycCnt[11]_net_1\, N_404, 
        \PrState_ns_0_0_0_a3_0_0[4]\, N_186_1, 
        CycCntlde_0_0_a3_0_0, \PrState[0]_net_1\, 
        \PrState[3]_net_1\, Phase2Cnt_n15_0_0_0_a3_0, 
        \Phase2Cnt[15]_net_1\, Phase2Cnt_n15_0_0_0_a3_0_0, N_144, 
        \PrState_ns_i_a3_i_0_o2_1[3]\, \Phase2Cnt[2]_net_1\, 
        \Phase2Cnt[3]_net_1\, \PrState_ns_i_a3_i_0_o2_0[3]\, 
        \Phase2Cnt[8]_net_1\, Phase2Cnt_n14_0_0_0_a3_0, 
        \Phase2Cnt[14]_net_1\, Phase2Cnt_n14_0_0_0_a3_0_0, 
        Phase2Cnt_n13_0_0_0_a3_0, \Phase2Cnt[13]_net_1\, 
        Phase2Cnt_n13_0_0_0_a3_0_0, Phase2Cnt_n12_0_0_0_a3_0, 
        \Phase2Cnt[12]_net_1\, Phase2Cnt_n12_0_0_0_a3_0_0, 
        Phase2Cnt_n11_0_0_0_a3_0, \Phase2Cnt[11]_net_1\, 
        Phase2Cnt_n11_0_0_0_a3_0_0, Phase2Cnt_n10_0_0_0_a3_0, 
        \Phase2Cnt[10]_net_1\, Phase2Cnt_n10_0_0_0_a3_0_0, 
        Phase2Cnt_n9_0_0_0_a3_0, \Phase2Cnt[9]_net_1\, 
        \PrState[1]_net_1\, Phase2Cnt_n9_0_0_0_a3_0_0, 
        Phase2Cnt_n6_0_i_0_0, N_169, \Phase2Cnt[6]_net_1\, 
        Phase2Cnt_n4_0_i_0_0, N_133, N_111, 
        \PrState_ns_i_a3_i_0_a3_0_0[3]\, N_242_9, 
        Phase2Cnt_n3_0_i_0_0, \PrState_ns_i_0_0_a3_1[0]\, 
        \PrState[4]_net_1\, \PrState_ns_i_0_0_a3_0[0]\, 
        \PrState_ns_0_i_0_a3_1_10_5[2]\, 
        \PrState_ns_0_i_0_a3_1_10_3[2]\, \Phase1Cnt[6]_net_1\, 
        \Phase1Cnt[5]_net_1\, \PrState_ns_0_i_0_a3_1_10_4[2]\, 
        \Phase1Cnt[4]_net_1\, \Phase1Cnt[3]_net_1\, 
        \PrState_ns_0_i_0_a3_1_10_1[2]\, \Phase1Cnt[0]_net_1\, 
        \Phase1Cnt[7]_net_1\, \Phase1Cnt[1]_net_1\, 
        \Phase1Cnt[2]_net_1\, \PrState_ns_0_i_0_a3_1_9_1[2]\, 
        \Phase1Cnt[9]_net_1\, \Phase1Cnt[10]_net_1\, 
        \PrState_ns_0_i_0_a3_1_9_0[2]\, \Phase1Cnt[11]_net_1\, 
        \Phase1Cnt[8]_net_1\, N_28, \Phase2Cnt[0]_net_1\, 
        \Phase2Cnt[1]_net_1\, N_32, N_188, N_167, N_34, 
        \Phase2Cnt[4]_net_1\, N_36, N_190, N_38, N_114, N_40, 
        N_192, N_172, N_42, N_171, N_193, N_20, N_141, N_433, 
        N_24, \CycCnt[8]_net_1\, N_145, N_162, N_402, N_207, 
        N_204, N_203, N_147, N_200, N_199, N_139, N_196, N_195, 
        \Phase2Cnt[7]_net_1\, N_22_i_0, \CycCnt[7]_net_1\, N_18, 
        \CycCnt[5]_net_1\, N_136, N_16, \CycCnt[4]_net_1\, N_135, 
        N_14, \CycCnt[3]_net_1\, N_119, N_12, \CycCnt[2]_net_1\, 
        N_113, N_10, \CycCnt[0]_net_1\, \CycCnt[1]_net_1\, N_227, 
        N_242_10, N_243, N_23, N_233, N_398, N_25, N_27, N_400, 
        N_21, N_146, N_19, N_231, N_17, N_140, N_15, N_137, 
        N_13_i_0, Phase2Cnt_n0, \Phase2Cnt[5]_net_1\, 
        \CycCnt[6]_net_1\, CycCnte, N_30, N_174_i_i_0, 
        Phase2Cnt_n9, Phase2Cnt_n10, Phase2Cnt_n11, N_179, 
        Phase2Cnt_n12, Phase2Cnt_n13, N_177, Phase2Cnt_n14, 
        Phase2Cnt_n15, N_175, \PrState_RNO_7[3]\, 
        \PrState_RNO_0[3]_net_1\, CycCnt_n9, \CycCnt[9]_net_1\, 
        N_397, CycCnt_n11, N_401, \DelayCnt[0]_net_1\, 
        \CycCnt[10]_net_1\, CycCnt_n10, CycCnt_n0, Phase1Cnt_n0, 
        \PrState_RNO_4[2]\, \PrState_ns[4]\, N_185, 
        \PrState_RNO_2[4]\, Phase1Cnt_n9, N_403, Phase1Cnt_n10, 
        N_407, N_173, Phase1Cnt_n11, \lvdsFifoRowRdOut\, \GND\, 
        \VCC\, GND_0, VCC_0 : std_logic;

begin 

    lvdsFifoRowRdOut <= \lvdsFifoRowRdOut\;

    \PrState[2]\ : DFN1C0
      port map(D => \PrState_RNO_4[2]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \PrState[2]_net_1\);
    
    \Phase2Cnt_RNO[7]\ : NOR3A
      port map(A => \PrState[1]_net_1\, B => N_192, C => N_172, Y
         => N_40);
    
    \Phase2Cnt_RNINV5B[2]\ : NOR2B
      port map(A => \Phase2Cnt[3]_net_1\, B => 
        \Phase2Cnt[2]_net_1\, Y => N_133);
    
    \PrState_RNO[0]\ : AO1B
      port map(A => \PrState_ns_0_0_0_a3_0_0[4]\, B => N_162, C
         => N_185, Y => \PrState_ns[4]\);
    
    \PrState_RNIVSEC3[4]\ : AO1
      port map(A => CycCntlde_0_0_a3_0_0, B => N_162, C => 
        \PrState[4]_net_1\, Y => CycCnte);
    
    \PrState_RNO_1[4]\ : OR2
      port map(A => \PrState[1]_net_1\, B => \PrState[4]_net_1\, 
        Y => \PrState_ns_i_0_0_a3_1[0]\);
    
    \Phase2Cnt_RNIMD79[15]\ : OR2
      port map(A => \Phase2Cnt[8]_net_1\, B => 
        \Phase2Cnt[15]_net_1\, Y => \PrState_ns_i_a3_i_0_o2_0[3]\);
    
    \Phase2Cnt_RNO_1[9]\ : OR3B
      port map(A => N_114, B => \Phase2Cnt[7]_net_1\, C => 
        Phase2Cnt_n9_0_0_0_a3_0_0, Y => N_195);
    
    \Phase1Cnt[1]\ : DFN1C0
      port map(D => N_13_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[1]_net_1\);
    
    \Phase1Cnt_RNO[4]\ : NOR3A
      port map(A => \PrState[2]_net_1\, B => N_231, C => N_146, Y
         => N_19);
    
    \Phase2Cnt_RNO_1[10]\ : OAI1
      port map(A => N_139, B => N_144, C => 
        Phase2Cnt_n10_0_0_0_a3_0, Y => N_196);
    
    \DelayCnt[0]\ : DFN1C0
      port map(D => N_166, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \DelayCnt[0]_net_1\);
    
    WFO_RNI10K2 : INV
      port map(A => \lvdsFifoRowRdOut\, Y => lvdsFifoRowRdOut_i);
    
    \Phase2Cnt_RNO_0[2]\ : AX1E
      port map(A => \Phase2Cnt[0]_net_1\, B => 
        \Phase2Cnt[1]_net_1\, C => \Phase2Cnt[2]_net_1\, Y => 
        N_174_i_i_0);
    
    \Phase2Cnt_RNO_2[10]\ : NOR2B
      port map(A => \Phase2Cnt[10]_net_1\, B => 
        \PrState_0[1]_net_1\, Y => Phase2Cnt_n10_0_0_0_a3_0);
    
    \Phase1Cnt_RNITC571[6]\ : NOR3C
      port map(A => N_146, B => \Phase1Cnt[5]_net_1\, C => 
        \Phase1Cnt[6]_net_1\, Y => N_398);
    
    \CycCnt_RNIQ88U[3]\ : NOR2B
      port map(A => N_119, B => \CycCnt[3]_net_1\, Y => N_135);
    
    \CycCnt_RNI3BQ51[4]\ : NOR2B
      port map(A => N_135, B => \CycCnt[4]_net_1\, Y => N_136);
    
    \Phase2Cnt_RNIMSMD2[14]\ : NOR3B
      port map(A => N_402, B => \Phase2Cnt[14]_net_1\, C => 
        \PrState_ns_i_a3_i_0_o2_1[3]\, Y => N_162);
    
    \Phase1Cnt[5]\ : DFN1C0
      port map(D => N_21, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[5]_net_1\);
    
    \Phase2Cnt_RNO[0]\ : NOR2A
      port map(A => \PrState[1]_net_1\, B => \Phase2Cnt[0]_net_1\, 
        Y => Phase2Cnt_n0);
    
    \CycCnt_RNO[2]\ : XA1B
      port map(A => \CycCnt[2]_net_1\, B => N_113, C => 
        \PrState[4]_net_1\, Y => N_12);
    
    \PrState_RNO_1[2]\ : AO1A
      port map(A => N_242, B => \PrState[2]_net_1\, C => N_166, Y
         => \PrState_ns_0_i_0_a3_0[2]\);
    
    \Phase2Cnt[12]\ : DFN1C0
      port map(D => Phase2Cnt_n12, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \Phase2Cnt[12]_net_1\);
    
    \CycCnt[10]\ : DFN1E1C0
      port map(D => CycCnt_n10, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[10]_net_1\);
    
    \Phase2Cnt[0]\ : DFN1C0
      port map(D => Phase2Cnt_n0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \Phase2Cnt[0]_net_1\);
    
    \Phase2Cnt_RNO[14]\ : AO1B
      port map(A => Phase2Cnt_n14_0_0_0_a3_0_0, B => N_402, C => 
        N_204, Y => Phase2Cnt_n14);
    
    \Phase2Cnt_RNIG8EE1[11]\ : NOR3B
      port map(A => \Phase2Cnt[10]_net_1\, B => 
        \Phase2Cnt[11]_net_1\, C => N_139, Y => N_147);
    
    \Phase2Cnt[2]\ : DFN1C0
      port map(D => N_30, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase2Cnt[2]_net_1\);
    
    \CycCnt_RNIVMKB2[9]\ : OR2A
      port map(A => \CycCnt[9]_net_1\, B => N_397, Y => N_401);
    
    \PrState_RNO[2]\ : OA1
      port map(A => N_243, B => \PrState_ns_0_i_0_a3_0[2]\, C => 
        CMOS_DrvX_0_LVDSen_2, Y => \PrState_RNO_4[2]\);
    
    \PrState_RNO_1[0]\ : OR2B
      port map(A => \PrState[0]_net_1\, B => CMOS_DrvX_0_LVDSen_2, 
        Y => N_185);
    
    \Phase2Cnt_RNO_0[10]\ : OR3A
      port map(A => \PrState_0[1]_net_1\, B => N_144, C => 
        \Phase2Cnt[10]_net_1\, Y => Phase2Cnt_n10_0_0_0_a3_0_0);
    
    \Phase2Cnt[13]\ : DFN1C0
      port map(D => Phase2Cnt_n13, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \Phase2Cnt[13]_net_1\);
    
    \Phase1Cnt_RNO[11]\ : XA1A
      port map(A => \Phase1Cnt[11]_net_1\, B => N_173, C => 
        \PrState[2]_net_1\, Y => Phase1Cnt_n11);
    
    \PrState_RNIVDOD[1]\ : NOR2B
      port map(A => \PrState[1]_net_1\, B => CMOS_DrvX_0_LVDSen_2, 
        Y => N_186_1);
    
    \Phase2Cnt_RNO_0[4]\ : AO1B
      port map(A => N_133, B => N_111, C => \PrState[1]_net_1\, Y
         => Phase2Cnt_n4_0_i_0_0);
    
    \Phase2Cnt_RNIDDDK[2]\ : OR3
      port map(A => \Phase2Cnt[2]_net_1\, B => 
        \Phase2Cnt[3]_net_1\, C => \PrState_ns_i_a3_i_0_o2_0[3]\, 
        Y => \PrState_ns_i_a3_i_0_o2_1[3]\);
    
    \PrState[4]\ : DFN1P0
      port map(D => \PrState_RNO_2[4]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, PRE => PLL_Test1_0_SysRst_O, Q
         => \PrState[4]_net_1\);
    
    \Phase2Cnt_RNIGLOG[4]\ : NOR3C
      port map(A => \Phase2Cnt[0]_net_1\, B => 
        \Phase2Cnt[1]_net_1\, C => \Phase2Cnt[4]_net_1\, Y => 
        N_111);
    
    \Phase1Cnt_RNIBDOG[2]\ : NOR2A
      port map(A => \Phase1Cnt[2]_net_1\, B => N_137, Y => N_140);
    
    \CycCnt_RNO[8]\ : XA1C
      port map(A => \CycCnt[8]_net_1\, B => N_145, C => 
        \PrState[4]_net_1\, Y => N_24);
    
    \Phase2Cnt_RNO[2]\ : NOR2A
      port map(A => \PrState[1]_net_1\, B => N_174_i_i_0, Y => 
        N_30);
    
    \Phase1Cnt[11]\ : DFN1C0
      port map(D => Phase1Cnt_n11, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[11]_net_1\);
    
    \Phase1Cnt_RNO[9]\ : XA1A
      port map(A => \Phase1Cnt[9]_net_1\, B => N_403, C => 
        \PrState[2]_net_1\, Y => Phase1Cnt_n9);
    
    \Phase1Cnt_RNISKCI1[8]\ : OR2B
      port map(A => \Phase1Cnt[8]_net_1\, B => N_400, Y => N_403);
    
    \Phase1Cnt_RNIAVBM[4]\ : NOR3C
      port map(A => \Phase1Cnt[4]_net_1\, B => 
        \Phase1Cnt[3]_net_1\, C => 
        \PrState_ns_0_i_0_a3_1_10_1[2]\, Y => 
        \PrState_ns_0_i_0_a3_1_10_4[2]\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \Phase1Cnt_RNO[7]\ : XA1
      port map(A => N_398, B => \Phase1Cnt[7]_net_1\, C => 
        \PrState[2]_net_1\, Y => N_25);
    
    \Phase2Cnt_RNO_0[9]\ : NOR2B
      port map(A => \Phase2Cnt[9]_net_1\, B => \PrState[1]_net_1\, 
        Y => Phase2Cnt_n9_0_0_0_a3_0);
    
    \Phase2Cnt_RNILNLL1[13]\ : NOR3C
      port map(A => N_147, B => \Phase2Cnt[12]_net_1\, C => 
        \Phase2Cnt[13]_net_1\, Y => N_402);
    
    \Phase1Cnt_RNIHF5B[1]\ : OR2B
      port map(A => \Phase1Cnt[1]_net_1\, B => 
        \Phase1Cnt[0]_net_1\, Y => N_137);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    \Phase2Cnt_RNO[10]\ : OAI1
      port map(A => N_139, B => Phase2Cnt_n10_0_0_0_a3_0_0, C => 
        N_196, Y => Phase2Cnt_n10);
    
    \Phase1Cnt[0]\ : DFN1C0
      port map(D => Phase1Cnt_n0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[0]_net_1\);
    
    \CycCnt_RNO[7]\ : XA1C
      port map(A => \CycCnt[7]_net_1\, B => N_141, C => 
        \PrState[4]_net_1\, Y => N_22_i_0);
    
    \Phase1Cnt[2]\ : DFN1C0
      port map(D => N_15, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[2]_net_1\);
    
    \CycCnt_RNO[4]\ : XA1B
      port map(A => \CycCnt[4]_net_1\, B => N_135, C => 
        \PrState[4]_net_1\, Y => N_16);
    
    \Phase2Cnt[3]\ : DFN1C0
      port map(D => N_32, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase2Cnt[3]_net_1\);
    
    \Phase2Cnt[7]\ : DFN1C0
      port map(D => N_40, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase2Cnt[7]_net_1\);
    
    \CycCnt_RNO_0[6]\ : AOI1
      port map(A => N_136, B => \CycCnt[5]_net_1\, C => 
        \CycCnt[6]_net_1\, Y => N_433);
    
    \Phase2Cnt_RNO_1[13]\ : OR3B
      port map(A => N_147, B => \Phase2Cnt[12]_net_1\, C => N_144, 
        Y => N_177);
    
    \Phase2Cnt_RNO_0[5]\ : AOI1
      port map(A => N_133, B => N_111, C => \Phase2Cnt[5]_net_1\, 
        Y => N_190);
    
    \CycCnt_RNILA5G2[10]\ : OR2A
      port map(A => \CycCnt[10]_net_1\, B => N_401, Y => N_404);
    
    WFO : DFN1C0
      port map(D => \PrState[2]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \lvdsFifoRowRdOut\);
    
    \Phase2Cnt_RNO_2[13]\ : OR3B
      port map(A => N_147, B => \Phase2Cnt[12]_net_1\, C => 
        Phase2Cnt_n13_0_0_0_a3_0_0, Y => N_203);
    
    \Phase2Cnt_RNO_0[7]\ : AOI1
      port map(A => N_133, B => N_114, C => \Phase2Cnt[7]_net_1\, 
        Y => N_192);
    
    \Phase1Cnt_RNO_0[4]\ : AOI1
      port map(A => \Phase1Cnt[3]_net_1\, B => N_140, C => 
        \Phase1Cnt[4]_net_1\, Y => N_231);
    
    \Phase2Cnt[6]\ : DFN1C0
      port map(D => N_38, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase2Cnt[6]_net_1\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \Phase1Cnt_RNO[0]\ : NOR2A
      port map(A => \PrState[2]_net_1\, B => \Phase1Cnt[0]_net_1\, 
        Y => Phase1Cnt_n0);
    
    \CycCnt[6]\ : DFN1E1C0
      port map(D => N_20, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[6]_net_1\);
    
    \Phase2Cnt_RNIAFBM[1]\ : NOR3C
      port map(A => \Phase2Cnt[0]_net_1\, B => 
        \Phase2Cnt[1]_net_1\, C => N_133, Y => N_167);
    
    \Phase2Cnt[10]\ : DFN1C0
      port map(D => Phase2Cnt_n10, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \Phase2Cnt[10]_net_1\);
    
    \Phase2Cnt_RNIFP671[9]\ : OR3C
      port map(A => N_114, B => \Phase2Cnt[7]_net_1\, C => 
        \Phase2Cnt[9]_net_1\, Y => N_139);
    
    \Phase2Cnt_RNIDDVR[6]\ : NOR3C
      port map(A => N_111, B => \Phase2Cnt[5]_net_1\, C => 
        \Phase2Cnt[6]_net_1\, Y => N_114);
    
    \Phase1Cnt_RNISUOC1[7]\ : NOR2B
      port map(A => \Phase1Cnt[7]_net_1\, B => N_398, Y => N_400);
    
    \Phase2Cnt_RNO_3[13]\ : OR3A
      port map(A => \PrState_0[1]_net_1\, B => N_144, C => 
        \Phase2Cnt[13]_net_1\, Y => Phase2Cnt_n13_0_0_0_a3_0_0);
    
    \Phase2Cnt_RNO_1[12]\ : AO1C
      port map(A => N_144, B => N_147, C => 
        Phase2Cnt_n12_0_0_0_a3_0, Y => N_200);
    
    \Phase2Cnt_RNO_0[13]\ : NOR2B
      port map(A => \Phase2Cnt[13]_net_1\, B => 
        \PrState_0[1]_net_1\, Y => Phase2Cnt_n13_0_0_0_a3_0);
    
    \Phase1Cnt[3]\ : DFN1C0
      port map(D => N_17, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[3]_net_1\);
    
    \Phase2Cnt_RNO_2[12]\ : NOR2B
      port map(A => \Phase2Cnt[12]_net_1\, B => 
        \PrState_0[1]_net_1\, Y => Phase2Cnt_n12_0_0_0_a3_0);
    
    \PrState[1]\ : DFN1C0
      port map(D => N_8, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \PrState[1]_net_1\);
    
    \Phase2Cnt[14]\ : DFN1C0
      port map(D => Phase2Cnt_n14, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \Phase2Cnt[14]_net_1\);
    
    \Phase1Cnt[7]\ : DFN1C0
      port map(D => N_25, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[7]_net_1\);
    
    \Phase2Cnt_RNO[15]\ : AO1B
      port map(A => Phase2Cnt_n15_0_0_0_a3_0, B => N_175, C => 
        N_207, Y => Phase2Cnt_n15);
    
    \Phase1Cnt_RNO[2]\ : XA1A
      port map(A => N_137, B => \Phase1Cnt[2]_net_1\, C => 
        \PrState[2]_net_1\, Y => N_15);
    
    \CycCnt[3]\ : DFN1E1C0
      port map(D => N_14, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[3]_net_1\);
    
    \PrState_RNO_0[0]\ : NOR3A
      port map(A => N_186_1, B => \CycCnt[11]_net_1\, C => N_404, 
        Y => \PrState_ns_0_0_0_a3_0_0[4]\);
    
    \PrState_RNO_0[4]\ : OR3
      port map(A => \PrState[0]_net_1\, B => \PrState[3]_net_1\, 
        C => \PrState[2]_net_1\, Y => \PrState_ns_i_0_0_a3_0[0]\);
    
    \Phase2Cnt_RNO_1[3]\ : OAI1
      port map(A => \Phase2Cnt[2]_net_1\, B => 
        \Phase2Cnt[3]_net_1\, C => \PrState[1]_net_1\, Y => 
        Phase2Cnt_n3_0_i_0_0);
    
    \Phase2Cnt_RNO_1[11]\ : OR3A
      port map(A => \Phase2Cnt[10]_net_1\, B => N_139, C => N_144, 
        Y => N_179);
    
    \DelayCnt_RNIEL39[0]\ : NOR2A
      port map(A => \PrState[3]_net_1\, B => \DelayCnt[0]_net_1\, 
        Y => N_166);
    
    \Phase2Cnt_RNO_2[11]\ : OR3B
      port map(A => \Phase2Cnt[10]_net_1\, B => 
        Phase2Cnt_n11_0_0_0_a3_0_0, C => N_139, Y => N_199);
    
    \Phase2Cnt_RNO_0[6]\ : OAI1
      port map(A => N_169, B => \Phase2Cnt[6]_net_1\, C => 
        \PrState[1]_net_1\, Y => Phase2Cnt_n6_0_i_0_0);
    
    \Phase1Cnt[6]\ : DFN1C0
      port map(D => N_23, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[6]_net_1\);
    
    \Phase2Cnt[8]\ : DFN1C0
      port map(D => N_42, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase2Cnt[8]_net_1\);
    
    \Phase2Cnt[15]\ : DFN1C0
      port map(D => Phase2Cnt_n15, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \Phase2Cnt[15]_net_1\);
    
    \Phase2Cnt_RNO_1[14]\ : AO1C
      port map(A => N_144, B => N_402, C => 
        Phase2Cnt_n14_0_0_0_a3_0, Y => N_204);
    
    \PrState_RNIRF0D2[2]\ : OR3C
      port map(A => \PrState_ns_i_a3_i_0_a3_0_0[3]\, B => 
        N_242_10, C => CMOS_DrvX_0_LVDSen_1, Y => N_227);
    
    \Phase2Cnt_RNO_2[14]\ : NOR2B
      port map(A => \Phase2Cnt[14]_net_1\, B => 
        \PrState_0[1]_net_1\, Y => Phase2Cnt_n14_0_0_0_a3_0);
    
    \Phase2Cnt_RNI4VOC1[7]\ : NOR3C
      port map(A => N_114, B => \Phase2Cnt[7]_net_1\, C => N_133, 
        Y => N_172);
    
    \Phase2Cnt_RNO[5]\ : NOR3A
      port map(A => \PrState[1]_net_1\, B => N_190, C => N_169, Y
         => N_36);
    
    \Phase2Cnt_RNO_0[12]\ : NOR3A
      port map(A => \PrState_0[1]_net_1\, B => N_144, C => 
        \Phase2Cnt[12]_net_1\, Y => Phase2Cnt_n12_0_0_0_a3_0_0);
    
    \CycCnt_RNIOFUK1[6]\ : OR3C
      port map(A => \CycCnt[5]_net_1\, B => N_136, C => 
        \CycCnt[6]_net_1\, Y => N_141);
    
    \CycCnt[0]\ : DFN1E1C0
      port map(D => CycCnt_n0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[0]_net_1\);
    
    \Phase2Cnt_RNO_3[11]\ : NOR3A
      port map(A => \PrState_0[1]_net_1\, B => N_144, C => 
        \Phase2Cnt[11]_net_1\, Y => Phase2Cnt_n11_0_0_0_a3_0_0);
    
    \CycCnt[8]\ : DFN1E1C0
      port map(D => N_24, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[8]_net_1\);
    
    \Phase2Cnt_RNO[8]\ : NOR3A
      port map(A => \PrState[1]_net_1\, B => N_171, C => N_193, Y
         => N_42);
    
    \PrState[3]\ : DFN1C0
      port map(D => \PrState_RNO_7[3]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \PrState[3]_net_1\);
    
    \Phase2Cnt_RNO_0[11]\ : NOR2B
      port map(A => \Phase2Cnt[11]_net_1\, B => 
        \PrState_0[1]_net_1\, Y => Phase2Cnt_n11_0_0_0_a3_0);
    
    \Phase1Cnt_RNIGH79[10]\ : NOR2B
      port map(A => \Phase1Cnt[9]_net_1\, B => 
        \Phase1Cnt[10]_net_1\, Y => 
        \PrState_ns_0_i_0_a3_1_9_1[2]\);
    
    \CycCnt_RNI4IGS1[7]\ : OR2A
      port map(A => \CycCnt[7]_net_1\, B => N_141, Y => N_145);
    
    \PrState[0]\ : DFN1C0
      port map(D => \PrState_ns[4]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \PrState[0]_net_1\);
    
    \Phase2Cnt_RNO_2[9]\ : OR3A
      port map(A => \PrState[1]_net_1\, B => N_144, C => 
        \Phase2Cnt[9]_net_1\, Y => Phase2Cnt_n9_0_0_0_a3_0_0);
    
    \PrState_RNI2U4Q[2]\ : NOR2B
      port map(A => \PrState[2]_net_1\, B => N_242_9, Y => 
        \PrState_ns_i_a3_i_0_a3_0_0[3]\);
    
    \Phase2Cnt_RNO[3]\ : NOR3
      port map(A => N_188, B => Phase2Cnt_n3_0_i_0_0, C => N_167, 
        Y => N_32);
    
    \CycCnt_RNO[1]\ : XA1B
      port map(A => \CycCnt[0]_net_1\, B => \CycCnt[1]_net_1\, C
         => \PrState[4]_net_1\, Y => N_10);
    
    \Phase2Cnt_RNO_0[14]\ : NOR3A
      port map(A => \PrState_0[1]_net_1\, B => N_144, C => 
        \Phase2Cnt[14]_net_1\, Y => Phase2Cnt_n14_0_0_0_a3_0_0);
    
    \Phase1Cnt[8]\ : DFN1C0
      port map(D => N_27, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[8]_net_1\);
    
    \Phase1Cnt_RNI0VEI[10]\ : NOR2B
      port map(A => \PrState_ns_0_i_0_a3_1_9_1[2]\, B => 
        \PrState_ns_0_i_0_a3_1_9_0[2]\, Y => N_242_9);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    \Phase1Cnt_RNI2LUR[4]\ : NOR3C
      port map(A => N_140, B => \Phase1Cnt[3]_net_1\, C => 
        \Phase1Cnt[4]_net_1\, Y => N_146);
    
    \Phase2Cnt_RNI5VH11[5]\ : NOR3C
      port map(A => N_111, B => \Phase2Cnt[5]_net_1\, C => N_133, 
        Y => N_169);
    
    \Phase1Cnt_RNIN76B[7]\ : NOR2A
      port map(A => \Phase1Cnt[0]_net_1\, B => 
        \Phase1Cnt[7]_net_1\, Y => 
        \PrState_ns_0_i_0_a3_1_10_3[2]\);
    
    \PrState_RNO_0[2]\ : NOR2A
      port map(A => N_162, B => \PrState_ns_0_i_0_a3_0_0[2]\, Y
         => N_243);
    
    \Phase1Cnt_RNO_0[6]\ : AOI1
      port map(A => \Phase1Cnt[5]_net_1\, B => N_146, C => 
        \Phase1Cnt[6]_net_1\, Y => N_233);
    
    \Phase2Cnt_RNO[6]\ : AOI1
      port map(A => N_133, B => N_114, C => Phase2Cnt_n6_0_i_0_0, 
        Y => N_38);
    
    \PrState_RNO_3[2]\ : NOR2B
      port map(A => N_242_10, B => N_242_9, Y => N_242);
    
    \Phase1Cnt_RNO_0[11]\ : OR2A
      port map(A => \Phase1Cnt[10]_net_1\, B => N_407, Y => N_173);
    
    \Phase2Cnt_RNO_0[8]\ : NOR2
      port map(A => \Phase2Cnt[8]_net_1\, B => N_172, Y => N_193);
    
    \Phase1Cnt_RNIIVCM[6]\ : NOR3A
      port map(A => \PrState_ns_0_i_0_a3_1_10_3[2]\, B => 
        \Phase1Cnt[6]_net_1\, C => \Phase1Cnt[5]_net_1\, Y => 
        \PrState_ns_0_i_0_a3_1_10_5[2]\);
    
    \CycCnt[4]\ : DFN1E1C0
      port map(D => N_16, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[4]_net_1\);
    
    \Phase1Cnt_RNO[10]\ : XA1A
      port map(A => \Phase1Cnt[10]_net_1\, B => N_407, C => 
        \PrState[2]_net_1\, Y => Phase1Cnt_n10);
    
    \Phase2Cnt_RNIOLPG[8]\ : OR2B
      port map(A => \Phase2Cnt[8]_net_1\, B => N_133, Y => N_144);
    
    \Phase1Cnt_RNITE0O1[9]\ : OR2A
      port map(A => \Phase1Cnt[9]_net_1\, B => N_403, Y => N_407);
    
    \CycCnt_RNO[5]\ : XA1B
      port map(A => \CycCnt[5]_net_1\, B => N_136, C => 
        \PrState[4]_net_1\, Y => N_18);
    
    \PrState_RNO_2[2]\ : OAI1
      port map(A => \CycCnt[11]_net_1\, B => N_404, C => 
        \PrState_0[1]_net_1\, Y => \PrState_ns_0_i_0_a3_0_0[2]\);
    
    \Phase2Cnt_RNO[1]\ : XA1
      port map(A => \Phase2Cnt[0]_net_1\, B => 
        \Phase2Cnt[1]_net_1\, C => \PrState[1]_net_1\, Y => N_28);
    
    \Phase2Cnt_RNO_0[3]\ : AOI1
      port map(A => \Phase2Cnt[1]_net_1\, B => 
        \Phase2Cnt[0]_net_1\, C => \Phase2Cnt[3]_net_1\, Y => 
        N_188);
    
    \PrState_RNO[3]\ : OA1
      port map(A => \PrState_RNO_0[3]_net_1\, B => 
        \PrState[4]_net_1\, C => CMOS_DrvX_0_LVDSen_2, Y => 
        \PrState_RNO_7[3]\);
    
    \Phase1Cnt_RNISUOC1[4]\ : NOR2B
      port map(A => \PrState_ns_0_i_0_a3_1_10_5[2]\, B => 
        \PrState_ns_0_i_0_a3_1_10_4[2]\, Y => N_242_10);
    
    \PrState_0[1]\ : DFN1C0
      port map(D => N_8, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \PrState_0[1]_net_1\);
    
    \CycCnt_RNO[0]\ : NOR2
      port map(A => \PrState[4]_net_1\, B => \CycCnt[0]_net_1\, Y
         => CycCnt_n0);
    
    \Phase2Cnt[11]\ : DFN1C0
      port map(D => Phase2Cnt_n11, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \Phase2Cnt[11]_net_1\);
    
    \CycCnt[7]\ : DFN1E1C0
      port map(D => N_22_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[7]_net_1\);
    
    \Phase2Cnt_RNO[11]\ : AO1B
      port map(A => Phase2Cnt_n11_0_0_0_a3_0, B => N_179, C => 
        N_199, Y => Phase2Cnt_n11);
    
    \CycCnt_RNIB44F[1]\ : NOR2B
      port map(A => \CycCnt[1]_net_1\, B => \CycCnt[0]_net_1\, Y
         => N_113);
    
    \Phase2Cnt_RNO[4]\ : OA1B
      port map(A => N_167, B => \Phase2Cnt[4]_net_1\, C => 
        Phase2Cnt_n4_0_i_0_0, Y => N_34);
    
    \Phase1Cnt_RNO[5]\ : XA1
      port map(A => N_146, B => \Phase1Cnt[5]_net_1\, C => 
        \PrState[2]_net_1\, Y => N_21);
    
    \Phase2Cnt[4]\ : DFN1C0
      port map(D => N_34, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase2Cnt[4]_net_1\);
    
    \Phase1Cnt_RNIJN5B[1]\ : NOR2
      port map(A => \Phase1Cnt[1]_net_1\, B => 
        \Phase1Cnt[2]_net_1\, Y => 
        \PrState_ns_0_i_0_a3_1_10_1[2]\);
    
    \CycCnt[1]\ : DFN1E1C0
      port map(D => N_10, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[1]_net_1\);
    
    \Phase2Cnt[9]\ : DFN1C0
      port map(D => Phase2Cnt_n9, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \Phase2Cnt[9]_net_1\);
    
    \CycCnt_RNO[10]\ : XA1C
      port map(A => \CycCnt[10]_net_1\, B => N_401, C => 
        \PrState[4]_net_1\, Y => CycCnt_n10);
    
    \CycCnt[11]\ : DFN1E1C0
      port map(D => CycCnt_n11, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[11]_net_1\);
    
    \Phase1Cnt[10]\ : DFN1C0
      port map(D => Phase1Cnt_n10, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[10]_net_1\);
    
    \CycCnt_RNII6MM[2]\ : NOR2B
      port map(A => N_113, B => \CycCnt[2]_net_1\, Y => N_119);
    
    \Phase1Cnt_RNO[8]\ : XA1
      port map(A => N_400, B => \Phase1Cnt[8]_net_1\, C => 
        \PrState[2]_net_1\, Y => N_27);
    
    \CycCnt_RNO[9]\ : XA1C
      port map(A => \CycCnt[9]_net_1\, B => N_397, C => 
        \PrState[4]_net_1\, Y => CycCnt_n9);
    
    \PrState_RNI5P1N[0]\ : NOR3
      port map(A => \PrState[0]_net_1\, B => \PrState[3]_net_1\, 
        C => \PrState[2]_net_1\, Y => CycCntlde_0_0_a3_0_0);
    
    \PrState_RNIGQF85[1]\ : AO1C
      port map(A => N_162, B => N_186_1, C => N_227, Y => N_8);
    
    \Phase2Cnt_RNO_1[15]\ : OR3B
      port map(A => N_402, B => \Phase2Cnt[14]_net_1\, C => N_144, 
        Y => N_175);
    
    \Phase2Cnt_RNO_2[15]\ : OR3B
      port map(A => N_402, B => \Phase2Cnt[14]_net_1\, C => 
        Phase2Cnt_n15_0_0_0_a3_0_0, Y => N_207);
    
    \Phase1Cnt_RNO[3]\ : XA1
      port map(A => N_140, B => \Phase1Cnt[3]_net_1\, C => 
        \PrState[2]_net_1\, Y => N_17);
    
    \CycCnt_RNO[3]\ : XA1B
      port map(A => \CycCnt[3]_net_1\, B => N_119, C => 
        \PrState[4]_net_1\, Y => N_14);
    
    \Phase1Cnt_RNIGD79[11]\ : NOR2A
      port map(A => \Phase1Cnt[11]_net_1\, B => 
        \Phase1Cnt[8]_net_1\, Y => \PrState_ns_0_i_0_a3_1_9_0[2]\);
    
    \Phase2Cnt[1]\ : DFN1C0
      port map(D => N_28, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase2Cnt[1]_net_1\);
    
    \CycCnt_RNO[11]\ : XA1C
      port map(A => \CycCnt[11]_net_1\, B => N_404, C => 
        \PrState[4]_net_1\, Y => CycCnt_n11);
    
    \Phase1Cnt_RNO[6]\ : NOR3A
      port map(A => \PrState[2]_net_1\, B => N_233, C => N_398, Y
         => N_23);
    
    \Phase2Cnt_RNI5LCI1[7]\ : NOR3B
      port map(A => N_114, B => \Phase2Cnt[7]_net_1\, C => N_144, 
        Y => N_171);
    
    \CycCnt_RNO[6]\ : NOR3A
      port map(A => N_141, B => N_433, C => \PrState[4]_net_1\, Y
         => N_20);
    
    \Phase2Cnt_RNO_3[15]\ : OR3A
      port map(A => \PrState_0[1]_net_1\, B => N_144, C => 
        \Phase2Cnt[15]_net_1\, Y => Phase2Cnt_n15_0_0_0_a3_0_0);
    
    \Phase1Cnt[4]\ : DFN1C0
      port map(D => N_19, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[4]_net_1\);
    
    \PrState_RNO[4]\ : OA1B
      port map(A => \PrState_ns_i_0_0_a3_0[0]\, B => 
        \PrState_ns_i_0_0_a3_1[0]\, C => CMOS_DrvX_0_LVDSen_2, Y
         => \PrState_RNO_2[4]\);
    
    \CycCnt_RNIHK242[8]\ : OR2A
      port map(A => \CycCnt[8]_net_1\, B => N_145, Y => N_397);
    
    \Phase1Cnt[9]\ : DFN1C0
      port map(D => Phase1Cnt_n9, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[9]_net_1\);
    
    \Phase2Cnt_RNO[13]\ : AO1B
      port map(A => Phase2Cnt_n13_0_0_0_a3_0, B => N_177, C => 
        N_203, Y => Phase2Cnt_n13);
    
    \PrState_RNO_0[3]\ : NOR2B
      port map(A => \PrState[3]_net_1\, B => \DelayCnt[0]_net_1\, 
        Y => \PrState_RNO_0[3]_net_1\);
    
    \Phase1Cnt_RNO[1]\ : XA1
      port map(A => \Phase1Cnt[0]_net_1\, B => 
        \Phase1Cnt[1]_net_1\, C => \PrState[2]_net_1\, Y => 
        N_13_i_0);
    
    \Phase2Cnt_RNO_0[15]\ : NOR2B
      port map(A => \Phase2Cnt[15]_net_1\, B => 
        \PrState_0[1]_net_1\, Y => Phase2Cnt_n15_0_0_0_a3_0);
    
    \CycCnt[5]\ : DFN1E1C0
      port map(D => N_18, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[5]_net_1\);
    
    \Phase2Cnt_RNO[12]\ : AO1B
      port map(A => Phase2Cnt_n12_0_0_0_a3_0_0, B => N_147, C => 
        N_200, Y => Phase2Cnt_n12);
    
    \Phase2Cnt[5]\ : DFN1C0
      port map(D => N_36, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase2Cnt[5]_net_1\);
    
    \CycCnt[9]\ : DFN1E1C0
      port map(D => CycCnt_n9, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[9]_net_1\);
    
    \CycCnt[2]\ : DFN1E1C0
      port map(D => N_12, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[2]_net_1\);
    
    \Phase2Cnt_RNO[9]\ : AO1C
      port map(A => N_171, B => Phase2Cnt_n9_0_0_0_a3_0, C => 
        N_195, Y => Phase2Cnt_n9);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3;
use proasic3.all;

entity WaveGenSingleZ14 is

    port( PrState_2               : in    std_logic;
          PrState_0               : in    std_logic_vector(4 to 4);
          PLL_Test1_0_SysRst_O    : in    std_logic;
          PLL_Test1_0_Sys_66M_Clk : in    std_logic;
          latch4acc_0_sqmuxa      : out   std_logic;
          FifoRowRdOut_1          : in    std_logic;
          FifoRowRdOut_0          : in    std_logic;
          latch4acc_0_sqmuxa_0    : out   std_logic;
          CMOS_DrvX_0_SDramEn_0   : in    std_logic;
          latch4acc_0_sqmuxa_1    : out   std_logic
        );

end WaveGenSingleZ14;

architecture DEF_ARCH of WaveGenSingleZ14 is 

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AOI1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component XA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OAI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal Data2accEn, \PrState_ns_i_0_1[2]\, N_65, 
        \PrState[2]_net_1\, \PrState_ns_i_0_0[2]\, 
        \PrState_ns_i_0_a5_0_0[2]\, \PrState_i[3]\, 
        \PrState_ns_i_0_a5_0[2]\, \Phase1Cnt_i[0]\, 
        \PrState_i[1]\, N_145_i_0, N_196, N_147_i_0, N_201, N_202, 
        N_34_i_0, \CycCnt[8]_net_1\, N_61, N_32_i_0, 
        \CycCnt[7]_net_1\, N_60, N_30, \CycCnt[6]_net_1\, N_59, 
        N_28, \CycCnt[5]_net_1\, N_41, N_26, \CycCnt[4]_net_1\, 
        N_39, N_24, \CycCnt[3]_net_1\, N_38, N_22, 
        \CycCnt[2]_net_1\, N_194, N_20, CycCnt_c0, 
        \CycCnt[1]_net_1\, N_64, \Phase2Cnt[1]_net_1\, N_192_i, 
        N_4, N_6, N_8, N_188_i, N_10, \DelayCnt[1]_net_1\, 
        N_143_i_0, CycCnte, N_63, \CycCnt[9]_net_1\, N_62, 
        CycCnt_n9, CycCnt_n0, \GND\, \VCC\, GND_0, VCC_0
         : std_logic;

begin 


    WFO : DFN1C0
      port map(D => \PrState[2]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => Data2accEn);
    
    \PrState[2]\ : DFN1C0
      port map(D => N_145_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \PrState[2]_net_1\);
    
    \PrState_RNO_3[2]\ : AOI1B
      port map(A => \PrState_ns_i_0_a5_0_0[2]\, B => 
        \PrState_i[3]\, C => FifoRowRdOut_0, Y => 
        \PrState_ns_i_0_0[2]\);
    
    \CycCnt_RNIEM53[2]\ : NOR2B
      port map(A => N_194, B => \CycCnt[2]_net_1\, Y => N_38);
    
    \CycCnt_RNI7G95[4]\ : NOR2B
      port map(A => N_39, B => \CycCnt[4]_net_1\, Y => N_41);
    
    \CycCnt[9]\ : DFN1E1C0
      port map(D => CycCnt_n9, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[9]_net_1\);
    
    \CycCnt_RNO[7]\ : XA1C
      port map(A => \CycCnt[7]_net_1\, B => N_60, C => 
        PrState_0(4), Y => N_32_i_0);
    
    WFO_RNI3R58_1 : NOR2B
      port map(A => Data2accEn, B => CMOS_DrvX_0_SDramEn_0, Y => 
        latch4acc_0_sqmuxa);
    
    \PrState_RNO_4[2]\ : NOR2B
      port map(A => \Phase1Cnt_i[0]\, B => \PrState_i[1]\, Y => 
        \PrState_ns_i_0_a5_0_0[2]\);
    
    \DelayCnt_RNO[1]\ : XA1B
      port map(A => \DelayCnt[1]_net_1\, B => N_188_i, C => 
        \PrState_i[3]\, Y => N_10);
    
    \Phase2Cnt_RNIS882[1]\ : NOR3A
      port map(A => \Phase2Cnt[1]_net_1\, B => N_192_i, C => 
        \PrState_i[1]\, Y => N_63);
    
    \Phase2Cnt_RNO[1]\ : XA1B
      port map(A => N_192_i, B => \Phase2Cnt[1]_net_1\, C => 
        \PrState_i[1]\, Y => N_6);
    
    \CycCnt[8]\ : DFN1E1C0
      port map(D => N_34_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[8]_net_1\);
    
    \CycCnt[5]\ : DFN1E1C0
      port map(D => N_28, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[5]_net_1\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \CycCnt_RNO[4]\ : XA1B
      port map(A => \CycCnt[4]_net_1\, B => N_39, C => PrState_2, 
        Y => N_26);
    
    \CycCnt[0]\ : DFN1E1C0
      port map(D => CycCnt_n0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => CycCnte, Q => CycCnt_c0);
    
    \CycCnt_RNO[9]\ : XA1C
      port map(A => \CycCnt[9]_net_1\, B => N_62, C => PrState_2, 
        Y => CycCnt_n9);
    
    \PrState[1]\ : DFN1P0
      port map(D => N_147_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        PRE => PLL_Test1_0_SysRst_O, Q => \PrState_i[1]\);
    
    \CycCnt_RNO[6]\ : XA1B
      port map(A => \CycCnt[6]_net_1\, B => N_59, C => 
        PrState_0(4), Y => N_30);
    
    \CycCnt_RNI5DB6[5]\ : NOR2B
      port map(A => N_41, B => \CycCnt[5]_net_1\, Y => N_59);
    
    \PrState_RNO_0[2]\ : NOR2A
      port map(A => \PrState_i[3]\, B => \PrState[2]_net_1\, Y
         => \PrState_ns_i_0_a5_0[2]\);
    
    \CycCnt[2]\ : DFN1E1C0
      port map(D => N_22, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[2]_net_1\);
    
    \CycCnt_RNO[3]\ : XA1B
      port map(A => \CycCnt[3]_net_1\, B => N_38, C => PrState_2, 
        Y => N_24);
    
    \CycCnt_RNO[2]\ : XA1B
      port map(A => \CycCnt[2]_net_1\, B => N_194, C => PrState_2, 
        Y => N_22);
    
    \PrState_RNO[2]\ : AOI1B
      port map(A => \PrState_ns_i_0_a5_0[2]\, B => N_196, C => 
        \PrState_ns_i_0_1[2]\, Y => N_145_i_0);
    
    \CycCnt_RNO[0]\ : NOR2
      port map(A => PrState_2, B => CycCnt_c0, Y => CycCnt_n0);
    
    \Phase2Cnt_RNIQ9F3[1]\ : OR2
      port map(A => PrState_2, B => N_63, Y => CycCnte);
    
    \CycCnt_RNIAJ74[3]\ : NOR2B
      port map(A => N_38, B => \CycCnt[3]_net_1\, Y => N_39);
    
    \CycCnt[6]\ : DFN1E1C0
      port map(D => N_30, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[6]_net_1\);
    
    \PrState_RNO_0[1]\ : OR2B
      port map(A => \PrState_i[1]\, B => N_64, Y => N_201);
    
    \Phase1Cnt[0]\ : DFN1P0
      port map(D => N_64, CLK => PLL_Test1_0_Sys_66M_Clk, PRE => 
        PLL_Test1_0_SysRst_O, Q => \Phase1Cnt_i[0]\);
    
    \DelayCnt[1]\ : DFN1C0
      port map(D => N_10, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \DelayCnt[1]_net_1\);
    
    \CycCnt[3]\ : DFN1E1C0
      port map(D => N_24, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[3]_net_1\);
    
    \Phase2Cnt_RNO[0]\ : NOR2
      port map(A => \PrState_i[1]\, B => N_192_i, Y => N_4);
    
    \PrState_RNO[1]\ : OR3C
      port map(A => N_201, B => N_202, C => FifoRowRdOut_0, Y => 
        N_147_i_0);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \CycCnt_RNO[1]\ : XA1B
      port map(A => CycCnt_c0, B => \CycCnt[1]_net_1\, C => 
        PrState_2, Y => N_20);
    
    \CycCnt[1]\ : DFN1E1C0
      port map(D => N_20, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[1]_net_1\);
    
    \Phase1Cnt_RNI87O1[0]\ : OR2B
      port map(A => \PrState[2]_net_1\, B => \Phase1Cnt_i[0]\, Y
         => N_64);
    
    \CycCnt_RNIJP32[1]\ : NOR2B
      port map(A => \CycCnt[1]_net_1\, B => CycCnt_c0, Y => N_194);
    
    WFO_RNI3R58_0 : NOR2B
      port map(A => Data2accEn, B => CMOS_DrvX_0_SDramEn_0, Y => 
        latch4acc_0_sqmuxa_0);
    
    \Phase2Cnt[1]\ : DFN1C0
      port map(D => N_6, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase2Cnt[1]_net_1\);
    
    \DelayCnt[0]\ : DFN1C0
      port map(D => N_8, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => N_188_i);
    
    \CycCnt_RNI4AD7[6]\ : OR2B
      port map(A => N_59, B => \CycCnt[6]_net_1\, Y => N_60);
    
    \CycCnt_RNI54H9[8]\ : OR2A
      port map(A => \CycCnt[8]_net_1\, B => N_61, Y => N_62);
    
    \CycCnt[4]\ : DFN1E1C0
      port map(D => N_26, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[4]_net_1\);
    
    \PrState_RNO[3]\ : OAI1
      port map(A => N_65, B => PrState_2, C => FifoRowRdOut_1, Y
         => N_143_i_0);
    
    WFO_RNI3R58 : NOR2B
      port map(A => Data2accEn, B => CMOS_DrvX_0_SDramEn_0, Y => 
        latch4acc_0_sqmuxa_1);
    
    \CycCnt[7]\ : DFN1E1C0
      port map(D => N_32_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[7]_net_1\);
    
    \PrState[3]\ : DFN1P0
      port map(D => N_143_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        PRE => PLL_Test1_0_SysRst_O, Q => \PrState_i[3]\);
    
    \PrState_RNO_1[2]\ : OAI1
      port map(A => \CycCnt[9]_net_1\, B => N_62, C => N_63, Y
         => N_196);
    
    \CycCnt_RNI47F8[7]\ : OR2A
      port map(A => \CycCnt[7]_net_1\, B => N_60, Y => N_61);
    
    \CycCnt_RNO[5]\ : XA1B
      port map(A => \CycCnt[5]_net_1\, B => N_41, C => 
        PrState_0(4), Y => N_28);
    
    \DelayCnt_RNI2UF9[1]\ : OA1C
      port map(A => \DelayCnt[1]_net_1\, B => N_188_i, C => 
        \PrState_i[3]\, Y => N_65);
    
    \CycCnt_RNO[8]\ : XA1C
      port map(A => \CycCnt[8]_net_1\, B => N_61, C => 
        PrState_0(4), Y => N_34_i_0);
    
    \PrState_RNO_2[2]\ : OA1A
      port map(A => N_65, B => \PrState[2]_net_1\, C => 
        \PrState_ns_i_0_0[2]\, Y => \PrState_ns_i_0_1[2]\);
    
    \PrState_RNO_1[1]\ : OR3A
      port map(A => \Phase2Cnt[1]_net_1\, B => N_192_i, C => 
        \PrState[2]_net_1\, Y => N_202);
    
    \Phase2Cnt[0]\ : DFN1C0
      port map(D => N_4, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => N_192_i);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    \DelayCnt_RNO[0]\ : NOR2
      port map(A => \PrState_i[3]\, B => N_188_i, Y => N_8);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3;
use proasic3.all;

entity WaveGenSingleZ8 is

    port( lvdsFifoRowRdOut_i      : in    std_logic;
          Main_ctl4SD_0_ByteRdEn  : out   std_logic;
          PLL_Test1_0_SysRst_O    : in    std_logic;
          PLL_Test1_0_Sys_66M_Clk : in    std_logic;
          lvdsFifoRowRdOut        : in    std_logic
        );

end WaveGenSingleZ8;

architecture DEF_ARCH of WaveGenSingleZ8 is 

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component OAI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1E
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \PrState_ns_0_0_0[2]\, \PrState_ns_0_0_a2_1_3[2]\, 
        N_50, N_67, \PrState_ns_0_0_a2_0[2]\, \PrState[2]_net_1\, 
        \PrState_ns_0_0_a2_0_1[3]\, N_70_1, \PrState_ns_0_i_0[1]\, 
        \PrState[3]_net_1\, \PrState[4]_net_1\, 
        \PrState_ns_0_0_a2_1_1[2]\, \PrState_ns_0_0_a2_1_0[2]\, 
        \DelayCnt[3]_net_1\, \DelayCnt[4]_net_1\, 
        \DelayCnt[2]_net_1\, \PrState_ns_0_i_a2_0_2[1]\, 
        \PrState_ns_0_i_a2_0_1[1]\, \CycCnt_5_i_o2_0[0]\, 
        \PrState[0]_net_1\, \Phase2Cnt[0]_net_1\, N_26_i_0, 
        \Phase1Cnt[0]_net_1\, \Phase1Cnt[1]_net_1\, N_28_i_0, 
        N_44, \Phase1Cnt[4]_net_1\, N_30, N_45, 
        \Phase1Cnt[5]_net_1\, N_53, \CycCnt[0]_net_1\, N_69, 
        \PrState[1]_net_1\, N_10, \PrState_ns[2]\, N_111, N_58, 
        N_36, N_49, \Phase1Cnt_RNO_0[8]_net_1\, N_34, N_47, 
        \Phase1Cnt[7]_net_1\, N_32, N_46, \Phase1Cnt[6]_net_1\, 
        N_21, N_51, N_19, N_17, \DelayCnt[0]_net_1\, 
        \DelayCnt[1]_net_1\, Phase1Cnt_n0, Phase1Cnt_n10, 
        \Phase1Cnt[10]_net_1\, N_52, Phase1Cnt_n11, 
        \Phase1Cnt[11]_net_1\, N_55, \Phase1Cnt[3]_net_1\, N_187, 
        \Phase1Cnt_RNO_2[2]\, N_11_i, N_7, \Phase1Cnt[2]_net_1\, 
        N_117, N_61, N_54, \Phase1Cnt[9]_net_1\, 
        \Phase1Cnt[8]_net_1\, N_23, N_14, \PrState_ns[3]\, N_6, 
        Phase1Cnt_n9, DelayCnt_n0, \GND\, \VCC\, GND_0, VCC_0
         : std_logic;

begin 


    WFO : DFN1C0
      port map(D => \PrState[2]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => Main_ctl4SD_0_ByteRdEn);
    
    \PrState[2]\ : DFN1C0
      port map(D => \PrState_ns[2]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \PrState[2]_net_1\);
    
    \PrState_RNO_3[2]\ : NOR3C
      port map(A => \PrState_ns_0_0_a2_1_1[2]\, B => 
        \PrState_ns_0_0_a2_1_0[2]\, C => lvdsFifoRowRdOut, Y => 
        \PrState_ns_0_0_a2_1_3[2]\);
    
    \Phase1Cnt[4]\ : DFN1C0
      port map(D => N_28_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[4]_net_1\);
    
    \DelayCnt_RNO_0[4]\ : NOR2B
      port map(A => N_51, B => \DelayCnt[3]_net_1\, Y => N_54);
    
    \Phase1Cnt_RNO[4]\ : XA1
      port map(A => N_44, B => \Phase1Cnt[4]_net_1\, C => 
        \PrState[2]_net_1\, Y => N_28_i_0);
    
    \PrState_RNO_0[0]\ : NOR2A
      port map(A => N_53, B => \CycCnt[0]_net_1\, Y => N_61);
    
    \Phase1Cnt[1]\ : DFN1C0
      port map(D => N_26_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[1]_net_1\);
    
    \Phase1Cnt[11]\ : DFN1C0
      port map(D => Phase1Cnt_n11, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[11]_net_1\);
    
    \PrState_RNO_4[2]\ : OR3C
      port map(A => N_53, B => \CycCnt[0]_net_1\, C => 
        lvdsFifoRowRdOut, Y => N_67);
    
    \DelayCnt_RNO[1]\ : XA1
      port map(A => \DelayCnt[0]_net_1\, B => \DelayCnt[1]_net_1\, 
        C => \PrState[3]_net_1\, Y => N_17);
    
    \Phase1Cnt[5]\ : DFN1C0
      port map(D => N_30, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[5]_net_1\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \Phase1Cnt_RNO[2]\ : NOR2A
      port map(A => \PrState[2]_net_1\, B => N_11_i, Y => 
        \Phase1Cnt_RNO_2[2]\);
    
    \CycCnt[0]\ : DFN1C0
      port map(D => N_6, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \CycCnt[0]_net_1\);
    
    \PrState_RNO_1[3]\ : OAI1
      port map(A => \PrState[3]_net_1\, B => \PrState[4]_net_1\, 
        C => lvdsFifoRowRdOut, Y => \PrState_ns_0_i_0[1]\);
    
    \Phase1Cnt_RNO[1]\ : XA1
      port map(A => \Phase1Cnt[0]_net_1\, B => 
        \Phase1Cnt[1]_net_1\, C => \PrState[2]_net_1\, Y => 
        N_26_i_0);
    
    \Phase1Cnt_RNIG3T11[6]\ : NOR2B
      port map(A => \Phase1Cnt[6]_net_1\, B => N_46, Y => N_47);
    
    \PrState[1]\ : DFN1C0
      port map(D => \PrState_ns[3]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \PrState[1]_net_1\);
    
    \DelayCnt_RNO[4]\ : XA1
      port map(A => \DelayCnt[4]_net_1\, B => N_54, C => 
        \PrState[3]_net_1\, Y => N_23);
    
    \PrState_RNIK1T4[1]\ : NOR2A
      port map(A => \PrState[1]_net_1\, B => \Phase2Cnt[0]_net_1\, 
        Y => N_53);
    
    \Phase1Cnt_RNO[6]\ : XA1
      port map(A => N_46, B => \Phase1Cnt[6]_net_1\, C => 
        \PrState[2]_net_1\, Y => N_32);
    
    \Phase1Cnt_RNI9NP[11]\ : NOR2B
      port map(A => \Phase1Cnt[11]_net_1\, B => 
        \Phase1Cnt[10]_net_1\, Y => N_70_1);
    
    \PrState_RNO_0[2]\ : NOR2B
      port map(A => \PrState[2]_net_1\, B => lvdsFifoRowRdOut, Y
         => \PrState_ns_0_0_a2_0[2]\);
    
    \PrState_RNO[2]\ : AO1B
      port map(A => \PrState_ns_0_0_a2_0[2]\, B => N_111, C => 
        \PrState_ns_0_0_0[2]\, Y => \PrState_ns[2]\);
    
    \Phase1Cnt_RNIF1GG1_0[9]\ : NOR2
      port map(A => \Phase1Cnt[9]_net_1\, B => N_49, Y => N_117);
    
    \CycCnt_RNO[0]\ : XA1B
      port map(A => \CycCnt[0]_net_1\, B => N_58, C => 
        \PrState[4]_net_1\, Y => N_6);
    
    \DelayCnt[2]\ : DFN1C0
      port map(D => N_19, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \DelayCnt[2]_net_1\);
    
    \PrState_RNO_2[3]\ : NOR2
      port map(A => \DelayCnt[2]_net_1\, B => \DelayCnt[3]_net_1\, 
        Y => \PrState_ns_0_i_a2_0_1[1]\);
    
    \PrState_RNO_0[1]\ : NOR3C
      port map(A => N_70_1, B => \PrState[2]_net_1\, C => 
        lvdsFifoRowRdOut, Y => \PrState_ns_0_0_a2_0_1[3]\);
    
    \Phase1Cnt_RNIA9GE[2]\ : NOR3C
      port map(A => \Phase1Cnt[0]_net_1\, B => 
        \Phase1Cnt[1]_net_1\, C => \Phase1Cnt[2]_net_1\, Y => 
        N_187);
    
    \Phase1Cnt[0]\ : DFN1C0
      port map(D => Phase1Cnt_n0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[0]_net_1\);
    
    \Phase1Cnt_RNO[8]\ : NOR3B
      port map(A => \PrState[2]_net_1\, B => N_49, C => 
        \Phase1Cnt_RNO_0[8]_net_1\, Y => N_36);
    
    \DelayCnt[1]\ : DFN1C0
      port map(D => N_17, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \DelayCnt[1]_net_1\);
    
    \PrState_RNO_0[3]\ : NOR3B
      port map(A => \DelayCnt[4]_net_1\, B => 
        \PrState_ns_0_i_a2_0_1[1]\, C => \PrState[4]_net_1\, Y
         => \PrState_ns_0_i_a2_0_2[1]\);
    
    \Phase1Cnt_RNO[10]\ : XA1A
      port map(A => \Phase1Cnt[10]_net_1\, B => N_52, C => 
        \PrState[2]_net_1\, Y => Phase1Cnt_n10);
    
    \DelayCnt[3]\ : DFN1C0
      port map(D => N_21, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \DelayCnt[3]_net_1\);
    
    \PrState_RNO[1]\ : AO1B
      port map(A => \PrState_ns_0_0_a2_0_1[3]\, B => N_117, C => 
        N_69, Y => \PrState_ns[3]\);
    
    \PrState[4]\ : DFN1P0
      port map(D => lvdsFifoRowRdOut_i, CLK => 
        PLL_Test1_0_Sys_66M_Clk, PRE => PLL_Test1_0_SysRst_O, Q
         => \PrState[4]_net_1\);
    
    \DelayCnt_RNI12LC[1]\ : NOR2B
      port map(A => \DelayCnt[1]_net_1\, B => \DelayCnt[0]_net_1\, 
        Y => N_50);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \Phase1Cnt_RNIP8KB1[8]\ : OR3C
      port map(A => N_47, B => \Phase1Cnt[7]_net_1\, C => 
        \Phase1Cnt[8]_net_1\, Y => N_49);
    
    \Phase1Cnt_RNO[0]\ : NOR2A
      port map(A => \PrState[2]_net_1\, B => \Phase1Cnt[0]_net_1\, 
        Y => Phase1Cnt_n0);
    
    \Phase1Cnt[10]\ : DFN1C0
      port map(D => Phase1Cnt_n10, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[10]_net_1\);
    
    \DelayCnt_RNO[2]\ : XA1
      port map(A => \DelayCnt[2]_net_1\, B => N_50, C => 
        \PrState[3]_net_1\, Y => N_19);
    
    \Phase1Cnt_RNIF1GG1[9]\ : OR2A
      port map(A => \Phase1Cnt[9]_net_1\, B => N_49, Y => N_52);
    
    \DelayCnt_RNI3JVI[2]\ : NOR2B
      port map(A => N_50, B => \DelayCnt[2]_net_1\, Y => N_51);
    
    \DelayCnt[4]\ : DFN1C0
      port map(D => N_23, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \DelayCnt[4]_net_1\);
    
    \DelayCnt_RNO[3]\ : XA1
      port map(A => \DelayCnt[3]_net_1\, B => N_51, C => 
        \PrState[3]_net_1\, Y => N_21);
    
    \DelayCnt[0]\ : DFN1C0
      port map(D => DelayCnt_n0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \DelayCnt[0]_net_1\);
    
    \PrState[0]\ : DFN1C0
      port map(D => N_14, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \PrState[0]_net_1\);
    
    \Phase1Cnt[6]\ : DFN1C0
      port map(D => N_32, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[6]_net_1\);
    
    \PrState_RNO_6[2]\ : NOR2A
      port map(A => \DelayCnt[4]_net_1\, B => \DelayCnt[2]_net_1\, 
        Y => \PrState_ns_0_0_a2_1_0[2]\);
    
    \Phase1Cnt_RNIQ9BJ[3]\ : NOR2B
      port map(A => \Phase1Cnt[3]_net_1\, B => N_187, Y => N_44);
    
    \PrState_RNO_5[2]\ : NOR2A
      port map(A => \PrState[3]_net_1\, B => \DelayCnt[3]_net_1\, 
        Y => \PrState_ns_0_0_a2_1_1[2]\);
    
    \Phase1Cnt_RNO_0[2]\ : AX1E
      port map(A => \Phase1Cnt[0]_net_1\, B => 
        \Phase1Cnt[1]_net_1\, C => \Phase1Cnt[2]_net_1\, Y => 
        N_11_i);
    
    \Phase1Cnt_RNO[7]\ : XA1
      port map(A => N_47, B => \Phase1Cnt[7]_net_1\, C => 
        \PrState[2]_net_1\, Y => N_34);
    
    \Phase1Cnt[7]\ : DFN1C0
      port map(D => N_34, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[7]_net_1\);
    
    \Phase1Cnt_RNO[9]\ : XA1A
      port map(A => N_49, B => \Phase1Cnt[9]_net_1\, C => 
        \PrState[2]_net_1\, Y => Phase1Cnt_n9);
    
    \PrState_RNO[3]\ : AOI1
      port map(A => \PrState_ns_0_i_a2_0_2[1]\, B => N_50, C => 
        \PrState_ns_0_i_0[1]\, Y => N_10);
    
    \Phase1Cnt_RNITM1T[5]\ : NOR2A
      port map(A => \Phase1Cnt[5]_net_1\, B => N_45, Y => N_46);
    
    \PrState[3]\ : DFN1C0
      port map(D => N_10, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \PrState[3]_net_1\);
    
    \Phase1Cnt_RNO[3]\ : XA1
      port map(A => N_187, B => \Phase1Cnt[3]_net_1\, C => 
        \PrState[2]_net_1\, Y => N_7);
    
    \Phase1Cnt_RNO_0[8]\ : AOI1
      port map(A => \Phase1Cnt[7]_net_1\, B => N_47, C => 
        \Phase1Cnt[8]_net_1\, Y => \Phase1Cnt_RNO_0[8]_net_1\);
    
    \Phase1Cnt[9]\ : DFN1C0
      port map(D => Phase1Cnt_n9, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[9]_net_1\);
    
    \CycCnt_RNO_1[0]\ : OR2
      port map(A => \PrState[0]_net_1\, B => \Phase2Cnt[0]_net_1\, 
        Y => \CycCnt_5_i_o2_0[0]\);
    
    \PrState_RNO_1[2]\ : OR2B
      port map(A => N_117, B => N_70_1, Y => N_111);
    
    \PrState_RNO[0]\ : OA1
      port map(A => N_61, B => \PrState[0]_net_1\, C => 
        lvdsFifoRowRdOut, Y => N_14);
    
    \Phase1Cnt_RNIBE6O[4]\ : OR2B
      port map(A => \Phase1Cnt[4]_net_1\, B => N_44, Y => N_45);
    
    \Phase1Cnt_RNO_0[11]\ : OR2A
      port map(A => \Phase1Cnt[10]_net_1\, B => N_52, Y => N_55);
    
    \Phase1Cnt[3]\ : DFN1C0
      port map(D => N_7, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[3]_net_1\);
    
    \Phase1Cnt_RNO[5]\ : XA1A
      port map(A => N_45, B => \Phase1Cnt[5]_net_1\, C => 
        \PrState[2]_net_1\, Y => N_30);
    
    \CycCnt_RNO_0[0]\ : NOR3
      port map(A => \CycCnt_5_i_o2_0[0]\, B => \PrState[3]_net_1\, 
        C => \PrState[2]_net_1\, Y => N_58);
    
    \Phase1Cnt_RNO[11]\ : XA1A
      port map(A => \Phase1Cnt[11]_net_1\, B => N_55, C => 
        \PrState[2]_net_1\, Y => Phase1Cnt_n11);
    
    \PrState_RNO_2[2]\ : AOI1B
      port map(A => \PrState_ns_0_0_a2_1_3[2]\, B => N_50, C => 
        N_67, Y => \PrState_ns_0_0_0[2]\);
    
    \PrState_RNO_1[1]\ : OR3C
      port map(A => \Phase2Cnt[0]_net_1\, B => \PrState[1]_net_1\, 
        C => lvdsFifoRowRdOut, Y => N_69);
    
    \Phase2Cnt[0]\ : DFN1C0
      port map(D => N_53, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase2Cnt[0]_net_1\);
    
    \Phase1Cnt[8]\ : DFN1C0
      port map(D => N_36, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[8]_net_1\);
    
    \Phase1Cnt[2]\ : DFN1C0
      port map(D => \Phase1Cnt_RNO_2[2]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \Phase1Cnt[2]_net_1\);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    \DelayCnt_RNO[0]\ : NOR2A
      port map(A => \PrState[3]_net_1\, B => \DelayCnt[0]_net_1\, 
        Y => DelayCnt_n0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3;
use proasic3.all;

entity WaveGenSingleZ12 is

    port( PrState_4               : out   std_logic;
          PrState_0               : out   std_logic_vector(4 to 4);
          latch_en                : out   std_logic;
          FifoRowRdOut            : in    std_logic;
          FifoRowRdOut_0          : in    std_logic;
          PLL_Test1_0_SysRst_O    : in    std_logic;
          FifoRowRdOut_i          : in    std_logic;
          PLL_Test1_0_Sys_66M_Clk : in    std_logic
        );

end WaveGenSingleZ12;

architecture DEF_ARCH of WaveGenSingleZ12 is 

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AOI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1E
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OAI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \PrState_ns_0_i_0[1]\, \PrState[3]_net_1\, 
        \PrState_0[4]_net_1\, \PrState_ns_0_i_a2_0_0_0[1]\, 
        \DelayCnt[1]_net_1\, \DelayCnt[2]_net_1\, 
        \DelayCnt[0]_net_1\, \CycCnt_5_i_o2_0[0]\, 
        \PrState[0]_net_1\, \Phase2Cnt[0]_net_1\, N_19_i_0, 
        \Phase1Cnt[0]_net_1\, \Phase1Cnt[1]_net_1\, 
        \PrState[2]_net_1\, N_21_i_0, N_39, \Phase1Cnt[2]_net_1\, 
        N_23, N_40, \Phase1Cnt[3]_net_1\, N_25, N_167, N_42, N_27, 
        \Phase1Cnt[5]_net_1\, N_29, N_169, N_44, N_31, 
        \Phase1Cnt[7]_net_1\, N_33, N_45, \Phase1Cnt[8]_net_1\, 
        N_8, N_64, \PrState[1]_net_1\, N_54, N_14, 
        \PrState_ns_0_0_a2_1_1[2]\, DelayCnt_n0, 
        \PrState_ns_0_0_0[2]\, \PrState_ns_0_0_a2_0_0[2]\, N_49, 
        \CycCnt[0]_net_1\, \PrState_ns[2]\, N_51, N_65_1, 
        Phase1Cnt_n0, \Phase1Cnt[4]_net_1\, \Phase1Cnt[6]_net_1\, 
        Phase1Cnt_n9, \Phase1Cnt[9]_net_1\, N_46, Phase1Cnt_n10, 
        \Phase1Cnt[10]_net_1\, N_47, N_48, 
        \PrState_RNO_0[0]_net_1\, N_55_i, \Phase1Cnt[11]_net_1\, 
        Phase1Cnt_n11, N_16, N_12_i_0, \PrState_ns[3]\, N_6, 
        \PrState[4]_net_1\, \GND\, \VCC\, GND_0, VCC_0
         : std_logic;

begin 

    PrState_4 <= \PrState[4]_net_1\;
    PrState_0(4) <= \PrState_0[4]_net_1\;

    WFO : DFN1C0
      port map(D => \PrState[2]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => latch_en);
    
    \PrState[2]\ : DFN1C0
      port map(D => \PrState_ns[2]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \PrState[2]_net_1\);
    
    \Phase1Cnt_RNO_0[6]\ : AOI1
      port map(A => \Phase1Cnt[5]_net_1\, B => N_42, C => 
        \Phase1Cnt[6]_net_1\, Y => N_169);
    
    \Phase1Cnt[4]\ : DFN1C0
      port map(D => N_25, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[4]_net_1\);
    
    \DelayCnt_RNO_0[2]\ : AX1E
      port map(A => \DelayCnt[0]_net_1\, B => \DelayCnt[1]_net_1\, 
        C => \DelayCnt[2]_net_1\, Y => N_55_i);
    
    \Phase1Cnt_RNO[4]\ : NOR3A
      port map(A => \PrState[2]_net_1\, B => N_167, C => N_42, Y
         => N_25);
    
    \Phase1Cnt_RNION4E[8]\ : OR2B
      port map(A => \Phase1Cnt[8]_net_1\, B => N_45, Y => N_46);
    
    \PrState_RNO_0[0]\ : NOR2A
      port map(A => N_49, B => \CycCnt[0]_net_1\, Y => 
        \PrState_RNO_0[0]_net_1\);
    
    \Phase1Cnt[1]\ : DFN1C0
      port map(D => N_19_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[1]_net_1\);
    
    \Phase1Cnt[11]\ : DFN1C0
      port map(D => Phase1Cnt_n11, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[11]_net_1\);
    
    \DelayCnt_RNO[1]\ : XA1
      port map(A => \DelayCnt[0]_net_1\, B => \DelayCnt[1]_net_1\, 
        C => \PrState[3]_net_1\, Y => N_14);
    
    \Phase1Cnt[5]\ : DFN1C0
      port map(D => N_27, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[5]_net_1\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \PrState_RNIF673[2]\ : NOR2B
      port map(A => \PrState[2]_net_1\, B => FifoRowRdOut, Y => 
        N_65_1);
    
    \Phase1Cnt_RNO[2]\ : XA1A
      port map(A => N_39, B => \Phase1Cnt[2]_net_1\, C => 
        \PrState[2]_net_1\, Y => N_21_i_0);
    
    \PrState_RNIAVQ2[1]\ : NOR2A
      port map(A => \PrState[1]_net_1\, B => \Phase2Cnt[0]_net_1\, 
        Y => N_49);
    
    \CycCnt[0]\ : DFN1C0
      port map(D => N_6, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \CycCnt[0]_net_1\);
    
    \PrState_RNO_1[3]\ : OAI1
      port map(A => \PrState[3]_net_1\, B => \PrState_0[4]_net_1\, 
        C => FifoRowRdOut_0, Y => \PrState_ns_0_i_0[1]\);
    
    \Phase1Cnt_RNO[1]\ : XA1
      port map(A => \Phase1Cnt[0]_net_1\, B => 
        \Phase1Cnt[1]_net_1\, C => \PrState[2]_net_1\, Y => 
        N_19_i_0);
    
    \PrState[1]\ : DFN1C0
      port map(D => \PrState_ns[3]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \PrState[1]_net_1\);
    
    \Phase1Cnt_RNIL1NF[9]\ : OR2A
      port map(A => \Phase1Cnt[9]_net_1\, B => N_46, Y => N_47);
    
    \Phase1Cnt_RNO[6]\ : NOR3A
      port map(A => \PrState[2]_net_1\, B => N_169, C => N_44, Y
         => N_29);
    
    \PrState_RNO_0[2]\ : AO1B
      port map(A => \PrState_ns_0_0_a2_1_1[2]\, B => 
        \PrState_ns_0_0_a2_0_0[2]\, C => FifoRowRdOut_0, Y => 
        \PrState_ns_0_0_0[2]\);
    
    \PrState_RNO[2]\ : AO1C
      port map(A => N_51, B => N_65_1, C => \PrState_ns_0_0_0[2]\, 
        Y => \PrState_ns[2]\);
    
    \CycCnt_RNO[0]\ : XA1B
      port map(A => \CycCnt[0]_net_1\, B => N_54, C => 
        \PrState[4]_net_1\, Y => N_6);
    
    \DelayCnt[2]\ : DFN1C0
      port map(D => N_16, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \DelayCnt[2]_net_1\);
    
    \Phase1Cnt_RNI0K0O[11]\ : NOR2
      port map(A => \Phase1Cnt[11]_net_1\, B => N_48, Y => N_51);
    
    \PrState_RNO_0[1]\ : OR3C
      port map(A => \Phase2Cnt[0]_net_1\, B => \PrState[1]_net_1\, 
        C => FifoRowRdOut_0, Y => N_64);
    
    \Phase1Cnt_RNIVSM4[2]\ : OR2A
      port map(A => \Phase1Cnt[2]_net_1\, B => N_39, Y => N_40);
    
    \Phase1Cnt[0]\ : DFN1C0
      port map(D => Phase1Cnt_n0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[0]_net_1\);
    
    \Phase1Cnt_RNO[8]\ : XA1
      port map(A => N_45, B => \Phase1Cnt[8]_net_1\, C => 
        \PrState[2]_net_1\, Y => N_33);
    
    \DelayCnt[1]\ : DFN1C0
      port map(D => N_14, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \DelayCnt[1]_net_1\);
    
    \PrState_RNO_0[3]\ : NOR3B
      port map(A => \DelayCnt[1]_net_1\, B => \DelayCnt[2]_net_1\, 
        C => \DelayCnt[0]_net_1\, Y => 
        \PrState_ns_0_i_a2_0_0_0[1]\);
    
    \Phase1Cnt_RNO_0[4]\ : OA1C
      port map(A => \Phase1Cnt[3]_net_1\, B => N_40, C => 
        \Phase1Cnt[4]_net_1\, Y => N_167);
    
    \Phase1Cnt_RNO[10]\ : XA1A
      port map(A => \Phase1Cnt[10]_net_1\, B => N_47, C => 
        \PrState[2]_net_1\, Y => Phase1Cnt_n10);
    
    \Phase1Cnt_RNISDIC[7]\ : NOR2B
      port map(A => \Phase1Cnt[7]_net_1\, B => N_44, Y => N_45);
    
    \PrState_RNO[1]\ : AO1B
      port map(A => N_65_1, B => N_51, C => N_64, Y => 
        \PrState_ns[3]\);
    
    \PrState[4]\ : DFN1P0
      port map(D => FifoRowRdOut_i, CLK => 
        PLL_Test1_0_Sys_66M_Clk, PRE => PLL_Test1_0_SysRst_O, Q
         => \PrState[4]_net_1\);
    
    \PrState_0[4]\ : DFN1P0
      port map(D => FifoRowRdOut_i, CLK => 
        PLL_Test1_0_Sys_66M_Clk, PRE => PLL_Test1_0_SysRst_O, Q
         => \PrState_0[4]_net_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \Phase1Cnt_RNO[0]\ : NOR2A
      port map(A => \PrState[2]_net_1\, B => \Phase1Cnt[0]_net_1\, 
        Y => Phase1Cnt_n0);
    
    \Phase1Cnt_RNIQORJ[10]\ : OR2A
      port map(A => \Phase1Cnt[10]_net_1\, B => N_47, Y => N_48);
    
    \Phase1Cnt[10]\ : DFN1C0
      port map(D => Phase1Cnt_n10, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[10]_net_1\);
    
    \DelayCnt_RNO[2]\ : NOR2A
      port map(A => \PrState[3]_net_1\, B => N_55_i, Y => N_16);
    
    \Phase1Cnt_RNI9J43[1]\ : OR2B
      port map(A => \Phase1Cnt[1]_net_1\, B => 
        \Phase1Cnt[0]_net_1\, Y => N_39);
    
    \DelayCnt[0]\ : DFN1C0
      port map(D => DelayCnt_n0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \DelayCnt[0]_net_1\);
    
    \PrState[0]\ : DFN1C0
      port map(D => N_12_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \PrState[0]_net_1\);
    
    \DelayCnt_RNIK5H2[0]\ : NOR2A
      port map(A => \PrState[3]_net_1\, B => \DelayCnt[0]_net_1\, 
        Y => DelayCnt_n0);
    
    \Phase1Cnt[6]\ : DFN1C0
      port map(D => N_29, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[6]_net_1\);
    
    \Phase1Cnt_RNO[7]\ : XA1
      port map(A => N_44, B => \Phase1Cnt[7]_net_1\, C => 
        \PrState[2]_net_1\, Y => N_31);
    
    \Phase1Cnt[7]\ : DFN1C0
      port map(D => N_31, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[7]_net_1\);
    
    \Phase1Cnt_RNO[9]\ : XA1A
      port map(A => \Phase1Cnt[9]_net_1\, B => N_46, C => 
        \PrState[2]_net_1\, Y => Phase1Cnt_n9);
    
    \Phase1Cnt_RNIEGR7[4]\ : NOR3B
      port map(A => \Phase1Cnt[3]_net_1\, B => 
        \Phase1Cnt[4]_net_1\, C => N_40, Y => N_42);
    
    \PrState_RNO[3]\ : OA1C
      port map(A => \PrState_ns_0_i_a2_0_0_0[1]\, B => 
        \PrState_0[4]_net_1\, C => \PrState_ns_0_i_0[1]\, Y => 
        N_8);
    
    \PrState[3]\ : DFN1C0
      port map(D => N_8, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \PrState[3]_net_1\);
    
    \Phase1Cnt_RNO[3]\ : XA1A
      port map(A => N_40, B => \Phase1Cnt[3]_net_1\, C => 
        \PrState[2]_net_1\, Y => N_23);
    
    \Phase1Cnt[9]\ : DFN1C0
      port map(D => Phase1Cnt_n9, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[9]_net_1\);
    
    \CycCnt_RNO_1[0]\ : OR2
      port map(A => \PrState[0]_net_1\, B => \Phase2Cnt[0]_net_1\, 
        Y => \CycCnt_5_i_o2_0[0]\);
    
    \PrState_RNO_1[2]\ : OR3C
      port map(A => \DelayCnt[1]_net_1\, B => \DelayCnt[2]_net_1\, 
        C => DelayCnt_n0, Y => \PrState_ns_0_0_a2_1_1[2]\);
    
    \PrState_RNO[0]\ : OA1
      port map(A => \PrState_RNO_0[0]_net_1\, B => 
        \PrState[0]_net_1\, C => FifoRowRdOut, Y => N_12_i_0);
    
    \Phase1Cnt_RNI140B[6]\ : NOR3C
      port map(A => N_42, B => \Phase1Cnt[5]_net_1\, C => 
        \Phase1Cnt[6]_net_1\, Y => N_44);
    
    \Phase1Cnt[3]\ : DFN1C0
      port map(D => N_23, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[3]_net_1\);
    
    \Phase1Cnt_RNO[5]\ : XA1
      port map(A => N_42, B => \Phase1Cnt[5]_net_1\, C => 
        \PrState[2]_net_1\, Y => N_27);
    
    \CycCnt_RNO_0[0]\ : NOR3
      port map(A => \CycCnt_5_i_o2_0[0]\, B => \PrState[3]_net_1\, 
        C => \PrState[2]_net_1\, Y => N_54);
    
    \Phase1Cnt_RNO[11]\ : XA1A
      port map(A => \Phase1Cnt[11]_net_1\, B => N_48, C => 
        \PrState[2]_net_1\, Y => Phase1Cnt_n11);
    
    \PrState_RNO_2[2]\ : OR2B
      port map(A => N_49, B => \CycCnt[0]_net_1\, Y => 
        \PrState_ns_0_0_a2_0_0[2]\);
    
    \Phase2Cnt[0]\ : DFN1C0
      port map(D => N_49, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase2Cnt[0]_net_1\);
    
    \Phase1Cnt[8]\ : DFN1C0
      port map(D => N_33, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[8]_net_1\);
    
    \Phase1Cnt[2]\ : DFN1C0
      port map(D => N_21_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[2]_net_1\);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3;
use proasic3.all;

entity WaveGenSingleZ16 is

    port( PrState_2               : in    std_logic;
          PrState_0               : in    std_logic_vector(4 to 4);
          PLL_Test1_0_SysRst_O    : in    std_logic;
          PLL_Test1_0_Sys_66M_Clk : in    std_logic;
          lvds_fifoRd             : in    std_logic;
          Main_ctl4SD_0_fifo_rd   : out   std_logic;
          FifoRowRdOut_1          : in    std_logic;
          FifoRowRdOut_0          : in    std_logic
        );

end WaveGenSingleZ16;

architecture DEF_ARCH of WaveGenSingleZ16 is 

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component XA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NOR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OAI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \PrState_ns_i_0_1[2]\, N_84, N_83, 
        \PrState_ns_i_0_a5_0[2]\, \PrState[3]_net_1\, 
        \PrState[2]_net_1\, N_141_i_0, N_189, N_143_i_0, N_194, 
        N_195, \Phase1Cnt_i[0]\, \PrState_i[1]\, N_32_i_0, 
        \CycCnt[8]_net_1\, N_59, N_30_i_0, \CycCnt[7]_net_1\, 
        N_58, N_28, N_78, N_26, \CycCnt[5]_net_1\, N_39, N_24, 
        \CycCnt[4]_net_1\, N_37, N_22, \CycCnt[3]_net_1\, N_36, 
        N_20, \CycCnt[2]_net_1\, N_186, N_18, CycCnt_c0, 
        \CycCnt[1]_net_1\, N_62, \Phase2Cnt[1]_net_1\, N_184_i, 
        N_187, N_4, N_6, N_8, \DelayCnt[0]_net_1\, N_139_i_0, 
        CycCnte, N_61, \CycCnt[9]_net_1\, N_60, \CycCnt[6]_net_1\, 
        CycCnt_n9, CycCnt_n0, interFifo_rd, \GND\, \VCC\, GND_0, 
        VCC_0 : std_logic;

begin 


    WFO : DFN1C0
      port map(D => \PrState[2]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => interFifo_rd);
    
    \PrState[2]\ : DFN1C0
      port map(D => N_141_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \PrState[2]_net_1\);
    
    \PrState_RNO_3[2]\ : OR3B
      port map(A => \Phase1Cnt_i[0]\, B => \PrState_i[1]\, C => 
        \PrState[3]_net_1\, Y => N_84);
    
    \CycCnt_RNO_0[6]\ : AOI1
      port map(A => N_39, B => \CycCnt[5]_net_1\, C => 
        \CycCnt[6]_net_1\, Y => N_78);
    
    \CycCnt[9]\ : DFN1E1C0
      port map(D => CycCnt_n9, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[9]_net_1\);
    
    \CycCnt_RNO[7]\ : XA1C
      port map(A => \CycCnt[7]_net_1\, B => N_58, C => 
        PrState_0(4), Y => N_30_i_0);
    
    \PrState_RNO_4[2]\ : OR2
      port map(A => \PrState[2]_net_1\, B => N_187, Y => N_83);
    
    WFO_RNIFNP3 : OR2
      port map(A => lvds_fifoRd, B => interFifo_rd, Y => 
        Main_ctl4SD_0_fifo_rd);
    
    \CycCnt_RNIOECB1[8]\ : OR2A
      port map(A => \CycCnt[8]_net_1\, B => N_59, Y => N_60);
    
    \Phase2Cnt_RNO[1]\ : XA1B
      port map(A => N_184_i, B => \Phase2Cnt[1]_net_1\, C => 
        \PrState_i[1]\, Y => N_6);
    
    \CycCnt[8]\ : DFN1E1C0
      port map(D => N_32_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[8]_net_1\);
    
    \CycCnt[5]\ : DFN1E1C0
      port map(D => N_26, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[5]_net_1\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \CycCnt_RNO[4]\ : XA1B
      port map(A => \CycCnt[4]_net_1\, B => N_37, C => 
        PrState_0(4), Y => N_24);
    
    \CycCnt[0]\ : DFN1E1C0
      port map(D => CycCnt_n0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => CycCnte, Q => CycCnt_c0);
    
    \CycCnt_RNO[9]\ : XA1C
      port map(A => \CycCnt[9]_net_1\, B => N_60, C => PrState_2, 
        Y => CycCnt_n9);
    
    \PrState[1]\ : DFN1P0
      port map(D => N_143_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        PRE => PLL_Test1_0_SysRst_O, Q => \PrState_i[1]\);
    
    \CycCnt_RNO[6]\ : NOR3A
      port map(A => N_58, B => N_78, C => PrState_0(4), Y => N_28);
    
    \PrState_RNO_0[2]\ : NOR2
      port map(A => \PrState[3]_net_1\, B => \PrState[2]_net_1\, 
        Y => \PrState_ns_i_0_a5_0[2]\);
    
    \CycCnt[2]\ : DFN1E1C0
      port map(D => N_20, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[2]_net_1\);
    
    \CycCnt_RNO[3]\ : XA1B
      port map(A => \CycCnt[3]_net_1\, B => N_36, C => 
        PrState_0(4), Y => N_22);
    
    \CycCnt_RNO[2]\ : XA1B
      port map(A => \CycCnt[2]_net_1\, B => N_186, C => 
        PrState_0(4), Y => N_20);
    
    \PrState_RNO[2]\ : AOI1B
      port map(A => \PrState_ns_i_0_a5_0[2]\, B => N_189, C => 
        \PrState_ns_i_0_1[2]\, Y => N_141_i_0);
    
    \CycCnt_RNO[0]\ : NOR2
      port map(A => PrState_2, B => CycCnt_c0, Y => CycCnt_n0);
    
    \CycCnt[6]\ : DFN1E1C0
      port map(D => N_28, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[6]_net_1\);
    
    \PrState_RNO_0[1]\ : OR2B
      port map(A => \PrState_i[1]\, B => N_62, Y => N_194);
    
    \Phase1Cnt[0]\ : DFN1P0
      port map(D => N_62, CLK => PLL_Test1_0_Sys_66M_Clk, PRE => 
        PLL_Test1_0_SysRst_O, Q => \Phase1Cnt_i[0]\);
    
    \CycCnt[3]\ : DFN1E1C0
      port map(D => N_22, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[3]_net_1\);
    
    \Phase2Cnt_RNO[0]\ : NOR2
      port map(A => \PrState_i[1]\, B => N_184_i, Y => N_4);
    
    \PrState_RNO[1]\ : OR3C
      port map(A => N_194, B => N_195, C => FifoRowRdOut_0, Y => 
        N_143_i_0);
    
    \DelayCnt_RNIISMB[0]\ : OR2B
      port map(A => \PrState[3]_net_1\, B => \DelayCnt[0]_net_1\, 
        Y => N_187);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \CycCnt_RNO[1]\ : XA1B
      port map(A => CycCnt_c0, B => \CycCnt[1]_net_1\, C => 
        PrState_0(4), Y => N_18);
    
    \CycCnt[1]\ : DFN1E1C0
      port map(D => N_18, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[1]_net_1\);
    
    \Phase2Cnt_RNIB7IK[1]\ : NOR3A
      port map(A => \Phase2Cnt[1]_net_1\, B => N_184_i, C => 
        \PrState_i[1]\, Y => N_61);
    
    \CycCnt_RNIE32O[4]\ : NOR2B
      port map(A => N_37, B => \CycCnt[4]_net_1\, Y => N_39);
    
    \CycCnt_RNISLH61[7]\ : OR2A
      port map(A => \CycCnt[7]_net_1\, B => N_58, Y => N_59);
    
    \Phase2Cnt[1]\ : DFN1C0
      port map(D => N_6, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase2Cnt[1]_net_1\);
    
    \DelayCnt[0]\ : DFN1C0
      port map(D => N_8, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \DelayCnt[0]_net_1\);
    
    \CycCnt_RNI9LJ9[1]\ : NOR2B
      port map(A => \CycCnt[1]_net_1\, B => CycCnt_c0, Y => N_186);
    
    \CycCnt_RNIMQ7J[3]\ : NOR2B
      port map(A => N_36, B => \CycCnt[3]_net_1\, Y => N_37);
    
    \CycCnt[4]\ : DFN1E1C0
      port map(D => N_24, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[4]_net_1\);
    
    \PrState_RNO[3]\ : OA1A
      port map(A => N_187, B => PrState_2, C => FifoRowRdOut_1, Y
         => N_139_i_0);
    
    \CycCnt[7]\ : DFN1E1C0
      port map(D => N_30_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[7]_net_1\);
    
    \PrState[3]\ : DFN1C0
      port map(D => N_139_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \PrState[3]_net_1\);
    
    \PrState_RNO_1[2]\ : OAI1
      port map(A => \CycCnt[9]_net_1\, B => N_60, C => N_61, Y
         => N_189);
    
    \Phase2Cnt_RNI98PL[1]\ : OR2
      port map(A => PrState_2, B => N_61, Y => CycCnte);
    
    \CycCnt_RNO[5]\ : XA1B
      port map(A => \CycCnt[5]_net_1\, B => N_39, C => 
        PrState_0(4), Y => N_26);
    
    \CycCnt_RNIVLDE[2]\ : NOR2B
      port map(A => N_186, B => \CycCnt[2]_net_1\, Y => N_36);
    
    \CycCnt_RNO[8]\ : XA1C
      port map(A => \CycCnt[8]_net_1\, B => N_59, C => 
        PrState_0(4), Y => N_32_i_0);
    
    \PrState_RNO_2[2]\ : NOR3C
      port map(A => N_84, B => N_83, C => FifoRowRdOut_0, Y => 
        \PrState_ns_i_0_1[2]\);
    
    \PrState_RNO_1[1]\ : OR3A
      port map(A => \Phase2Cnt[1]_net_1\, B => N_184_i, C => 
        \PrState[2]_net_1\, Y => N_195);
    
    \Phase2Cnt[0]\ : DFN1C0
      port map(D => N_4, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => N_184_i);
    
    \Phase1Cnt_RNI043D[0]\ : OR2B
      port map(A => \PrState[2]_net_1\, B => \Phase1Cnt_i[0]\, Y
         => N_62);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    \DelayCnt_RNO[0]\ : NOR2A
      port map(A => \PrState[3]_net_1\, B => \DelayCnt[0]_net_1\, 
        Y => N_8);
    
    \CycCnt_RNI11N11[6]\ : OR3C
      port map(A => \CycCnt[5]_net_1\, B => N_39, C => 
        \CycCnt[6]_net_1\, Y => N_58);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3;
use proasic3.all;

entity WaveGenSingleZ17 is

    port( FifoRowRdOut            : out   std_logic;
          CMOS_DrvX_0_SDramEn_0   : in    std_logic;
          FifoRowRdOut_i          : out   std_logic;
          FifoRowRdOut_0          : out   std_logic;
          FifoRowRdOut_1          : out   std_logic;
          PLL_Test1_0_SysRst_O    : in    std_logic;
          PLL_Test1_0_Sys_66M_Clk : in    std_logic;
          FifoRowRdOut_2          : out   std_logic
        );

end WaveGenSingleZ17;

architecture DEF_ARCH of WaveGenSingleZ17 is 

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OAI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component XA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component AO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1E
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component INV
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \PrState[2]_net_1\, \FifoRowRdOut_0\, 
        \PrState_ns_0_i_0_0[1]\, N_213, CycCntlde_0_0_a3_0, 
        \PrState[0]_net_1\, \PrState[3]_net_1\, 
        \PrState_ns_i_0_0_a3_0[0]\, \PrState[1]_net_1\, 
        \PrState_ns_i_a3_i_0_a2_8[3]\, \Phase1Cnt[0]_net_1\, 
        \PrState_ns_i_a3_i_0_a2_5[3]\, \Phase1Cnt[8]_net_1\, 
        \PrState_ns_i_a3_i_0_a2_7[3]\, 
        \PrState_ns_i_a3_i_0_a2_3[3]\, \Phase1Cnt[5]_net_1\, 
        \Phase1Cnt[4]_net_1\, \PrState_ns_i_a3_i_0_a2_6[3]\, 
        \Phase1Cnt[11]_net_1\, \Phase1Cnt[3]_net_1\, 
        \PrState_ns_i_a3_i_0_a2_1[3]\, \Phase1Cnt[9]_net_1\, 
        \Phase1Cnt[10]_net_1\, \Phase1Cnt[6]_net_1\, 
        \Phase1Cnt[7]_net_1\, \Phase1Cnt[1]_net_1\, 
        \Phase1Cnt[2]_net_1\, \PrState_ns_i_a3_i_0_o2_0[3]\, 
        \Phase2Cnt[4]_net_1\, \Phase2Cnt[0]_net_1\, N_152, N_218, 
        N_10, \DelayCnt[0]_net_1\, \DelayCnt[1]_net_1\, N_12, 
        \DelayCnt[2]_net_1\, N_120, N_14, \DelayCnt[3]_net_1\, 
        N_124, N_20, N_348, N_159, N_13, \Phase2Cnt[1]_net_1\, 
        N_276_i_0, N_277_i_0, N_105, \Phase1Cnt_RNO_1[3]\, N_107, 
        \Phase1Cnt_RNO[4]_net_1\, N_173, N_111, N_24, N_27, N_113, 
        \Phase1Cnt_RNO[7]_net_1\, N_115, \Phase1Cnt_RNO[8]_net_1\, 
        N_117, N_314, \CycCnt[4]_net_1\, N_108, 
        \PrState[4]_net_1\, N_315, \CycCnt[5]_net_1\, N_110, 
        N_318, \CycCnt[8]_net_1\, N_116, N_344, N_123, N_9, N_204, 
        N_7, N_153, N_154, N_164, N_199, 
        \PrState_ns_0_0_0_a3_0_0[4]\, N_200, N_317_i_0, 
        \CycCnt[7]_net_1\, N_114, N_316, N_190, N_313, 
        \CycCnt[3]_net_1\, N_106, N_8, \CycCnt[2]_net_1\, N_104, 
        N_312, \CycCnt[0]_net_1\, \CycCnt[1]_net_1\, N_18, N_346, 
        N_158, N_211, N_168, \CycCnt[11]_net_1\, N_343, 
        DelayCnt_n0, \Phase2Cnt[2]_net_1\, \Phase2Cnt[3]_net_1\, 
        Phase1Cnt_n0, Phase2Cnt_n0, \DelayCnt[4]_net_1\, N_16, 
        N_135_i, N_22, N_6, Phase1Cnt_n9, N_119, Phase1Cnt_n10, 
        N_125, Phase1Cnt_n11, N_347, CycCnt_n9, \CycCnt[9]_net_1\, 
        N_118, CycCnt_n10, \CycCnt[10]_net_1\, N_122, 
        \CycCnt[6]_net_1\, CycCnt_n11, \PrState_ns[4]\, 
        \PrState_RNO[4]_net_1\, CycCnte, CycCnt_n0, \GND\, \VCC\, 
        GND_0, VCC_0 : std_logic;

begin 

    FifoRowRdOut_0 <= \FifoRowRdOut_0\;

    \PrState[2]\ : DFN1C0
      port map(D => N_7, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \PrState[2]_net_1\);
    
    \Phase1Cnt_RNI670B[10]\ : NOR2
      port map(A => \Phase1Cnt[9]_net_1\, B => 
        \Phase1Cnt[10]_net_1\, Y => \PrState_ns_i_a3_i_0_a2_5[3]\);
    
    \CycCnt_RNIAC54[3]\ : NOR2B
      port map(A => N_106, B => \CycCnt[3]_net_1\, Y => N_108);
    
    \PrState_RNO[0]\ : AO1B
      port map(A => \PrState[0]_net_1\, B => 
        CMOS_DrvX_0_SDramEn_0, C => N_168, Y => \PrState_ns[4]\);
    
    \CycCnt_RNIFN65[4]\ : NOR2B
      port map(A => N_108, B => \CycCnt[4]_net_1\, Y => N_110);
    
    \Phase1Cnt_RNINNJC[1]\ : NOR2
      port map(A => \Phase1Cnt[1]_net_1\, B => 
        \Phase1Cnt[2]_net_1\, Y => \PrState_ns_i_a3_i_0_a2_1[3]\);
    
    \Phase1Cnt[1]\ : DFN1C0
      port map(D => N_276_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[1]_net_1\);
    
    \Phase1Cnt_RNO[4]\ : NOR3A
      port map(A => \PrState[2]_net_1\, B => N_173, C => N_111, Y
         => \Phase1Cnt_RNO[4]_net_1\);
    
    \PrState_RNI6V1D1[1]\ : NOR2A
      port map(A => N_344, B => N_211, Y => 
        \PrState_ns_0_0_0_a3_0_0[4]\);
    
    \DelayCnt[0]\ : DFN1C0
      port map(D => DelayCnt_n0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \DelayCnt[0]_net_1\);
    
    \Phase2Cnt_RNO_0[2]\ : AOI1
      port map(A => \Phase2Cnt[1]_net_1\, B => 
        \Phase2Cnt[0]_net_1\, C => \Phase2Cnt[2]_net_1\, Y => 
        N_158);
    
    \Phase1Cnt_RNIUF9P[4]\ : NOR3A
      port map(A => \PrState_ns_i_a3_i_0_a2_3[3]\, B => 
        \Phase1Cnt[5]_net_1\, C => \Phase1Cnt[4]_net_1\, Y => 
        \PrState_ns_i_a3_i_0_a2_7[3]\);
    
    \Phase1Cnt[5]\ : DFN1C0
      port map(D => N_24, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[5]_net_1\);
    
    \PrState_RNO[1]\ : OAI1
      port map(A => N_211, B => N_344, C => N_164, Y => N_6);
    
    \Phase2Cnt_RNO[0]\ : NOR2A
      port map(A => \PrState[1]_net_1\, B => \Phase2Cnt[0]_net_1\, 
        Y => Phase2Cnt_n0);
    
    \CycCnt_RNO[2]\ : XA1B
      port map(A => \CycCnt[2]_net_1\, B => N_104, C => 
        \PrState[4]_net_1\, Y => N_8);
    
    \PrState_RNO_1[2]\ : OR3B
      port map(A => \PrState[2]_net_1\, B => 
        CMOS_DrvX_0_SDramEn_0, C => N_218, Y => N_152);
    
    \Phase1Cnt_RNI2JKN[8]\ : NOR3B
      port map(A => \Phase1Cnt[0]_net_1\, B => 
        \PrState_ns_i_a3_i_0_a2_5[3]\, C => \Phase1Cnt[8]_net_1\, 
        Y => \PrState_ns_i_a3_i_0_a2_8[3]\);
    
    \CycCnt[10]\ : DFN1E1C0
      port map(D => CycCnt_n10, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[10]_net_1\);
    
    \Phase2Cnt[0]\ : DFN1C0
      port map(D => Phase2Cnt_n0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \Phase2Cnt[0]_net_1\);
    
    \PrState_RNIL9GD[1]\ : OR2B
      port map(A => \PrState[1]_net_1\, B => 
        CMOS_DrvX_0_SDramEn_0, Y => N_211);
    
    \Phase2Cnt[2]\ : DFN1C0
      port map(D => N_18, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase2Cnt[2]_net_1\);
    
    \PrState_RNO[2]\ : OR3C
      port map(A => N_153, B => N_152, C => N_154, Y => N_7);
    
    \Phase2Cnt_RNINPTI[3]\ : OR3C
      port map(A => \Phase2Cnt[1]_net_1\, B => 
        \Phase2Cnt[2]_net_1\, C => \Phase2Cnt[3]_net_1\, Y => 
        N_123);
    
    \Phase1Cnt_RNI10LC[6]\ : NOR2
      port map(A => \Phase1Cnt[6]_net_1\, B => 
        \Phase1Cnt[7]_net_1\, Y => \PrState_ns_i_a3_i_0_a2_3[3]\);
    
    \Phase1Cnt_RNO[11]\ : XA1A
      port map(A => \Phase1Cnt[11]_net_1\, B => N_347, C => 
        \PrState[2]_net_1\, Y => Phase1Cnt_n11);
    
    \Phase1Cnt_RNIELRO1[8]\ : OR2B
      port map(A => \Phase1Cnt[8]_net_1\, B => N_117, Y => N_119);
    
    \DelayCnt_RNO[3]\ : XA1
      port map(A => \DelayCnt[3]_net_1\, B => N_124, C => 
        \PrState[3]_net_1\, Y => N_14);
    
    \PrState[4]\ : DFN1P0
      port map(D => \PrState_RNO[4]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, PRE => PLL_Test1_0_SysRst_O, Q
         => \PrState[4]_net_1\);
    
    \CycCnt_RNO[8]\ : XA1C
      port map(A => \CycCnt[8]_net_1\, B => N_116, C => 
        \PrState[4]_net_1\, Y => N_318);
    
    \Phase2Cnt_RNO[2]\ : NOR3A
      port map(A => \PrState[1]_net_1\, B => N_346, C => N_158, Y
         => N_18);
    
    \Phase1Cnt_RNILFJC[1]\ : OR2B
      port map(A => \Phase1Cnt[1]_net_1\, B => 
        \Phase1Cnt[0]_net_1\, Y => N_105);
    
    \Phase1Cnt[11]\ : DFN1C0
      port map(D => Phase1Cnt_n11, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[11]_net_1\);
    
    \CycCnt_RNID4C9[8]\ : OR2A
      port map(A => \CycCnt[8]_net_1\, B => N_116, Y => N_118);
    
    \Phase1Cnt_RNO[9]\ : XA1A
      port map(A => \Phase1Cnt[9]_net_1\, B => N_119, C => 
        \PrState[2]_net_1\, Y => Phase1Cnt_n9);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \Phase1Cnt_RNO[7]\ : XA1
      port map(A => N_115, B => \Phase1Cnt[7]_net_1\, C => 
        \PrState[2]_net_1\, Y => \Phase1Cnt_RNO[7]_net_1\);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    \Phase1Cnt_RNIBD6C1[6]\ : NOR2B
      port map(A => \Phase1Cnt[6]_net_1\, B => N_113, Y => N_115);
    
    \PrState_RNIA90M1[4]\ : AO1
      port map(A => CycCntlde_0_0_a3_0, B => N_344, C => 
        \PrState[4]_net_1\, Y => CycCnte);
    
    \Phase1Cnt[0]\ : DFN1C0
      port map(D => Phase1Cnt_n0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[0]_net_1\);
    
    \CycCnt_RNO[7]\ : XA1C
      port map(A => \CycCnt[7]_net_1\, B => N_114, C => 
        \PrState[4]_net_1\, Y => N_317_i_0);
    
    \Phase1Cnt[2]\ : DFN1C0
      port map(D => N_277_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[2]_net_1\);
    
    \CycCnt_RNO[4]\ : XA1B
      port map(A => \CycCnt[4]_net_1\, B => N_108, C => 
        \PrState[4]_net_1\, Y => N_314);
    
    \DelayCnt[1]\ : DFN1C0
      port map(D => N_10, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \DelayCnt[1]_net_1\);
    
    \Phase2Cnt[3]\ : DFN1C0
      port map(D => N_20, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase2Cnt[3]_net_1\);
    
    \DelayCnt_RNIB8VN[4]\ : NOR3B
      port map(A => \DelayCnt[3]_net_1\, B => N_124, C => 
        \DelayCnt[4]_net_1\, Y => N_204);
    
    \CycCnt_RNO_0[6]\ : AOI1
      port map(A => N_110, B => \CycCnt[5]_net_1\, C => 
        \CycCnt[6]_net_1\, Y => N_190);
    
    WFO : DFN1C0
      port map(D => \PrState[2]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => FifoRowRdOut);
    
    \CycCnt_RNI4PA8[7]\ : OR2A
      port map(A => \CycCnt[7]_net_1\, B => N_114, Y => N_116);
    
    WFO_2 : DFN1C0
      port map(D => \PrState[2]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => FifoRowRdOut_2);
    
    \Phase1Cnt_RNO_0[4]\ : OA1C
      port map(A => \Phase1Cnt[3]_net_1\, B => N_107, C => 
        \Phase1Cnt[4]_net_1\, Y => N_173);
    
    \DelayCnt_RNO[4]\ : NOR2A
      port map(A => \PrState[3]_net_1\, B => N_135_i, Y => N_16);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \Phase1Cnt_RNO[0]\ : NOR2A
      port map(A => \PrState[2]_net_1\, B => \Phase1Cnt[0]_net_1\, 
        Y => Phase1Cnt_n0);
    
    \CycCnt[6]\ : DFN1E1C0
      port map(D => N_316, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[6]_net_1\);
    
    \Phase1Cnt_RNIO6JN[11]\ : NOR3C
      port map(A => \Phase1Cnt[11]_net_1\, B => 
        \Phase1Cnt[3]_net_1\, C => \PrState_ns_i_a3_i_0_a2_1[3]\, 
        Y => \PrState_ns_i_a3_i_0_a2_6[3]\);
    
    \DelayCnt_RNO[1]\ : XA1
      port map(A => \DelayCnt[0]_net_1\, B => \DelayCnt[1]_net_1\, 
        C => \PrState[3]_net_1\, Y => N_10);
    
    \DelayCnt[2]\ : DFN1C0
      port map(D => N_12, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \DelayCnt[2]_net_1\);
    
    \Phase1Cnt[3]\ : DFN1C0
      port map(D => \Phase1Cnt_RNO_1[3]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \Phase1Cnt[3]_net_1\);
    
    \PrState[1]\ : DFN1C0
      port map(D => N_6, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \PrState[1]_net_1\);
    
    \Phase1Cnt[7]\ : DFN1C0
      port map(D => \Phase1Cnt_RNO[7]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \Phase1Cnt[7]_net_1\);
    
    \Phase1Cnt_RNO[2]\ : XA1A
      port map(A => N_105, B => \Phase1Cnt[2]_net_1\, C => 
        \PrState[2]_net_1\, Y => N_277_i_0);
    
    \CycCnt[3]\ : DFN1E1C0
      port map(D => N_313, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[3]_net_1\);
    
    \PrState_RNO_0[0]\ : OR3A
      port map(A => \PrState_ns_0_0_0_a3_0_0[4]\, B => 
        \CycCnt[11]_net_1\, C => N_343, Y => N_168);
    
    \PrState_RNO_0[4]\ : OR3
      port map(A => \PrState[0]_net_1\, B => \PrState[2]_net_1\, 
        C => \PrState[1]_net_1\, Y => \PrState_ns_i_0_0_a3_0[0]\);
    
    \CycCnt_RNI9ORC[10]\ : OR2A
      port map(A => \CycCnt[10]_net_1\, B => N_122, Y => N_343);
    
    WFO_1 : DFN1C0
      port map(D => \PrState[2]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => FifoRowRdOut_1);
    
    \PrState_RNO_0[1]\ : OR3C
      port map(A => N_218, B => \PrState[2]_net_1\, C => 
        CMOS_DrvX_0_SDramEn_0, Y => N_164);
    
    \Phase1Cnt[6]\ : DFN1C0
      port map(D => N_27, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[6]_net_1\);
    
    \CycCnt_RNINFDA[9]\ : OR2A
      port map(A => \CycCnt[9]_net_1\, B => N_118, Y => N_122);
    
    \Phase1Cnt_RNIO9H82[11]\ : NOR3C
      port map(A => \PrState_ns_i_a3_i_0_a2_7[3]\, B => 
        \PrState_ns_i_a3_i_0_a2_6[3]\, C => 
        \PrState_ns_i_a3_i_0_a2_8[3]\, Y => N_218);
    
    \Phase1Cnt_RNIHDTI[2]\ : OR2A
      port map(A => \Phase1Cnt[2]_net_1\, B => N_105, Y => N_107);
    
    \CycCnt[0]\ : DFN1E1C0
      port map(D => CycCnt_n0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[0]_net_1\);
    
    \CycCnt[8]\ : DFN1E1C0
      port map(D => N_318, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[8]_net_1\);
    
    \PrState[3]\ : DFN1C0
      port map(D => N_9, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \PrState[3]_net_1\);
    
    \Phase1Cnt_RNICLHV[4]\ : NOR3B
      port map(A => \Phase1Cnt[3]_net_1\, B => 
        \Phase1Cnt[4]_net_1\, C => N_107, Y => N_111);
    
    \DelayCnt_RNO_0[4]\ : AX1E
      port map(A => \DelayCnt[3]_net_1\, B => N_124, C => 
        \DelayCnt[4]_net_1\, Y => N_135_i);
    
    \CycCnt_RNISD97[6]\ : OR3C
      port map(A => \CycCnt[5]_net_1\, B => N_110, C => 
        \CycCnt[6]_net_1\, Y => N_114);
    
    \PrState[0]\ : DFN1C0
      port map(D => \PrState_ns[4]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \PrState[0]_net_1\);
    
    \CycCnt_RNI6143[2]\ : NOR2B
      port map(A => N_104, B => \CycCnt[2]_net_1\, Y => N_106);
    
    \Phase2Cnt_RNO[3]\ : NOR3A
      port map(A => \PrState[1]_net_1\, B => N_348, C => N_159, Y
         => N_20);
    
    \DelayCnt[3]\ : DFN1C0
      port map(D => N_14, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \DelayCnt[3]_net_1\);
    
    \DelayCnt_RNIABCE[2]\ : NOR2B
      port map(A => N_120, B => \DelayCnt[2]_net_1\, Y => N_124);
    
    \CycCnt_RNO[1]\ : XA1B
      port map(A => \CycCnt[0]_net_1\, B => \CycCnt[1]_net_1\, C
         => \PrState[4]_net_1\, Y => N_312);
    
    \Phase1Cnt[8]\ : DFN1C0
      port map(D => \Phase1Cnt_RNO[8]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \Phase1Cnt[8]_net_1\);
    
    \Phase1Cnt_RNICVGI1[7]\ : NOR2B
      port map(A => \Phase1Cnt[7]_net_1\, B => N_115, Y => N_117);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    \PrState_RNIVJ7B[3]\ : OR2
      port map(A => \PrState[4]_net_1\, B => \PrState[3]_net_1\, 
        Y => N_213);
    
    \PrState_RNO_0[2]\ : OR3C
      port map(A => CMOS_DrvX_0_SDramEn_0, B => 
        \PrState[3]_net_1\, C => N_204, Y => N_153);
    
    \Phase2Cnt_RNIIF7P[0]\ : NOR2A
      port map(A => \Phase2Cnt[0]_net_1\, B => N_123, Y => N_348);
    
    \PrState_RNO_3[2]\ : OR3
      port map(A => \CycCnt[11]_net_1\, B => N_343, C => 
        \PrState[2]_net_1\, Y => N_199);
    
    \Phase1Cnt_RNO_0[11]\ : OR2A
      port map(A => \Phase1Cnt[10]_net_1\, B => N_125, Y => N_347);
    
    \CycCnt[4]\ : DFN1E1C0
      port map(D => N_314, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[4]_net_1\);
    
    \Phase1Cnt_RNO[10]\ : XA1A
      port map(A => \Phase1Cnt[10]_net_1\, B => N_125, C => 
        \PrState[2]_net_1\, Y => Phase1Cnt_n10);
    
    \CycCnt_RNO[5]\ : XA1B
      port map(A => \CycCnt[5]_net_1\, B => N_110, C => 
        \PrState[4]_net_1\, Y => N_315);
    
    \PrState_RNO_2[2]\ : OR3C
      port map(A => N_199, B => \PrState_ns_0_0_0_a3_0_0[4]\, C
         => N_200, Y => N_154);
    
    \Phase2Cnt_RNO[1]\ : XA1
      port map(A => \Phase2Cnt[0]_net_1\, B => 
        \Phase2Cnt[1]_net_1\, C => \PrState[1]_net_1\, Y => N_13);
    
    \Phase2Cnt_RNO_0[3]\ : NOR2
      port map(A => \Phase2Cnt[3]_net_1\, B => N_346, Y => N_159);
    
    \PrState_RNO[3]\ : OA1C
      port map(A => N_204, B => \PrState[4]_net_1\, C => 
        \PrState_ns_0_i_0_0[1]\, Y => N_9);
    
    \Phase2Cnt_RNIQRJC[4]\ : OR2
      port map(A => \Phase2Cnt[4]_net_1\, B => 
        \Phase2Cnt[0]_net_1\, Y => \PrState_ns_i_a3_i_0_o2_0[3]\);
    
    \CycCnt_RNO[0]\ : NOR2
      port map(A => \PrState[4]_net_1\, B => \CycCnt[0]_net_1\, Y
         => CycCnt_n0);
    
    WFO_0_RNI22P3 : INV
      port map(A => \FifoRowRdOut_0\, Y => FifoRowRdOut_i);
    
    \Phase1Cnt_RNIHF6V1[9]\ : OR2A
      port map(A => \Phase1Cnt[9]_net_1\, B => N_119, Y => N_125);
    
    \PrState_RNIPNQG[0]\ : NOR3
      port map(A => \PrState[0]_net_1\, B => \PrState[2]_net_1\, 
        C => \PrState[3]_net_1\, Y => CycCntlde_0_0_a3_0);
    
    \Phase1Cnt_RNIBVR51[5]\ : NOR2B
      port map(A => \Phase1Cnt[5]_net_1\, B => N_111, Y => N_113);
    
    \DelayCnt_RNO[2]\ : XA1
      port map(A => \DelayCnt[2]_net_1\, B => N_120, C => 
        \PrState[3]_net_1\, Y => N_12);
    
    \CycCnt[7]\ : DFN1E1C0
      port map(D => N_317_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[7]_net_1\);
    
    \Phase2Cnt_RNO[4]\ : XA1
      port map(A => N_348, B => \Phase2Cnt[4]_net_1\, C => 
        \PrState[1]_net_1\, Y => N_22);
    
    \Phase1Cnt_RNO[5]\ : XA1
      port map(A => N_111, B => \Phase1Cnt[5]_net_1\, C => 
        \PrState[2]_net_1\, Y => N_24);
    
    \Phase2Cnt_RNIHLHV[4]\ : NOR2
      port map(A => \PrState_ns_i_a3_i_0_o2_0[3]\, B => N_123, Y
         => N_344);
    
    \Phase2Cnt[4]\ : DFN1C0
      port map(D => N_22, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase2Cnt[4]_net_1\);
    
    \CycCnt[1]\ : DFN1E1C0
      port map(D => N_312, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[1]_net_1\);
    
    \CycCnt_RNO[10]\ : XA1C
      port map(A => \CycCnt[10]_net_1\, B => N_122, C => 
        \PrState[4]_net_1\, Y => CycCnt_n10);
    
    \CycCnt[11]\ : DFN1E1C0
      port map(D => CycCnt_n11, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[11]_net_1\);
    
    \Phase1Cnt[10]\ : DFN1C0
      port map(D => Phase1Cnt_n10, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[10]_net_1\);
    
    \Phase1Cnt_RNO[8]\ : XA1
      port map(A => N_117, B => \Phase1Cnt[8]_net_1\, C => 
        \PrState[2]_net_1\, Y => \Phase1Cnt_RNO[8]_net_1\);
    
    \CycCnt_RNO[9]\ : XA1C
      port map(A => \CycCnt[9]_net_1\, B => N_118, C => 
        \PrState[4]_net_1\, Y => CycCnt_n9);
    
    \DelayCnt_RNIRSI9[1]\ : NOR2B
      port map(A => \DelayCnt[1]_net_1\, B => \DelayCnt[0]_net_1\, 
        Y => N_120);
    
    \Phase1Cnt_RNO[3]\ : XA1A
      port map(A => N_107, B => \Phase1Cnt[3]_net_1\, C => 
        \PrState[2]_net_1\, Y => \Phase1Cnt_RNO_1[3]\);
    
    \CycCnt_RNO[3]\ : XA1B
      port map(A => \CycCnt[3]_net_1\, B => N_106, C => 
        \PrState[4]_net_1\, Y => N_313);
    
    \CycCnt_RNI3M22[1]\ : NOR2B
      port map(A => \CycCnt[1]_net_1\, B => \CycCnt[0]_net_1\, Y
         => N_104);
    
    \DelayCnt[4]\ : DFN1C0
      port map(D => N_16, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \DelayCnt[4]_net_1\);
    
    \DelayCnt_RNO[0]\ : NOR2A
      port map(A => \PrState[3]_net_1\, B => \DelayCnt[0]_net_1\, 
        Y => DelayCnt_n0);
    
    \Phase2Cnt[1]\ : DFN1C0
      port map(D => N_13, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase2Cnt[1]_net_1\);
    
    \CycCnt_RNO[11]\ : XA1C
      port map(A => \CycCnt[11]_net_1\, B => N_343, C => 
        \PrState[4]_net_1\, Y => CycCnt_n11);
    
    WFO_0 : DFN1C0
      port map(D => \PrState[2]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \FifoRowRdOut_0\);
    
    \Phase1Cnt_RNO[6]\ : XA1
      port map(A => N_113, B => \Phase1Cnt[6]_net_1\, C => 
        \PrState[2]_net_1\, Y => N_27);
    
    \CycCnt_RNO[6]\ : NOR3A
      port map(A => N_114, B => N_190, C => \PrState[4]_net_1\, Y
         => N_316);
    
    \Phase1Cnt[4]\ : DFN1C0
      port map(D => \Phase1Cnt_RNO[4]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \Phase1Cnt[4]_net_1\);
    
    \PrState_RNO[4]\ : OA1B
      port map(A => N_213, B => \PrState_ns_i_0_0_a3_0[0]\, C => 
        CMOS_DrvX_0_SDramEn_0, Y => \PrState_RNO[4]_net_1\);
    
    \PrState_RNO_4[2]\ : OR3A
      port map(A => N_218, B => \CycCnt[11]_net_1\, C => N_343, Y
         => N_200);
    
    \Phase1Cnt[9]\ : DFN1C0
      port map(D => Phase1Cnt_n9, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[9]_net_1\);
    
    \PrState_RNO_0[3]\ : OR2B
      port map(A => N_213, B => CMOS_DrvX_0_SDramEn_0, Y => 
        \PrState_ns_0_i_0_0[1]\);
    
    \Phase1Cnt_RNO[1]\ : XA1
      port map(A => \Phase1Cnt[0]_net_1\, B => 
        \Phase1Cnt[1]_net_1\, C => \PrState[2]_net_1\, Y => 
        N_276_i_0);
    
    \CycCnt[5]\ : DFN1E1C0
      port map(D => N_315, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[5]_net_1\);
    
    \Phase2Cnt_RNIKDTI[2]\ : NOR3C
      port map(A => \Phase2Cnt[1]_net_1\, B => 
        \Phase2Cnt[2]_net_1\, C => \Phase2Cnt[0]_net_1\, Y => 
        N_346);
    
    \CycCnt[9]\ : DFN1E1C0
      port map(D => CycCnt_n9, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[9]_net_1\);
    
    \CycCnt[2]\ : DFN1E1C0
      port map(D => N_8, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[2]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3;
use proasic3.all;

entity WaveGenSingleZ10 is

    port( lvds_fifoRd             : out   std_logic;
          PLL_Test1_0_SysRst_O    : in    std_logic;
          PLL_Test1_0_Sys_66M_Clk : in    std_logic;
          lvdsFifoRowRdOut        : in    std_logic
        );

end WaveGenSingleZ10;

architecture DEF_ARCH of WaveGenSingleZ10 is 

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1E
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component XA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component XAI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \PrState_ns_0_0_a2_0[2]\, N_78, N_67, 
        \PrState_ns_0_0_a2_0_0[4]\, \PrState_ns_0_i_0[1]\, N_150, 
        CycCntlde_0_a2_0_0, \PrState[0]_net_1\, 
        \PrState[2]_net_1\, \PrState[3]_net_1\, 
        \PrState_ns_i_0_a2_0[0]\, \PrState[1]_net_1\, 
        \PrState_ns_0_0_a2_0_2[2]\, \DelayCnt[0]_net_1\, 
        \DelayCnt[1]_net_1\, \PrState_ns_0_0_a2_0_0[2]\, 
        \DelayCnt[3]_net_1\, \PrState_ns_0_0_a2_0[3]\, 
        \PrState_ns_0_i_a2_1[1]\, \PrState[4]_net_1\, 
        \PrState_ns_0_i_a2_0_0[1]\, \PrState_ns_0_i_a2_0[1]\, 
        N_13, \CycCnt[0]_net_1\, \CycCnt[1]_net_1\, N_15, 
        \CycCnt[2]_net_1\, N_44, N_17, \CycCnt[3]_net_1\, N_177, 
        N_19, \CycCnt[4]_net_1\, N_46, N_21, \CycCnt[5]_net_1\, 
        N_47, N_23, N_68, N_192, N_25_i_0, \CycCnt[7]_net_1\, 
        N_27_i_0, \CycCnt[8]_net_1\, N_70, N_186_i, N_92, 
        \CycCnt[9]_net_1\, N_74, N_7, N_39, N_72, N_37, 
        \DelayCnt_i[2]\, N_69, N_35, N_33, N_116, N_117, N_31, 
        \Phase2Cnt[0]_net_1\, \Phase2Cnt[1]_net_1\, 
        \DelayCnt[4]_net_1\, CycCnt_n0, \CycCnt[6]_net_1\, 
        CycCnt_n9, CycCnte, N_73, N_79_i, \Phase2Cnt[2]_net_1\, 
        \Phase1Cnt[0]_net_1\, N_41, \PrState_ns[4]\, 
        \PrState_ns[3]\, N_90, \PrState_ns[2]\, N_129, 
        \PrState_RNO_3[4]\, NxState_0_sqmuxa, DelayCnt_n0, 
        Phase2Cnt_n0, \GND\, \VCC\, GND_0, VCC_0 : std_logic;

begin 


    WFO : DFN1C0
      port map(D => \PrState[2]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => lvds_fifoRd);
    
    \PrState[2]\ : DFN1C0
      port map(D => \PrState_ns[2]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \PrState[2]_net_1\);
    
    \PrState_RNO_3[2]\ : NOR2A
      port map(A => \PrState[3]_net_1\, B => \DelayCnt[3]_net_1\, 
        Y => \PrState_ns_0_0_a2_0_0[2]\);
    
    \CycCnt_RNI2E5L[3]\ : NOR2B
      port map(A => N_177, B => \CycCnt[3]_net_1\, Y => N_46);
    
    \DelayCnt_RNO_0[4]\ : AX1E
      port map(A => \DelayCnt[3]_net_1\, B => N_72, C => 
        \DelayCnt[4]_net_1\, Y => N_79_i);
    
    \DelayCnt_RNIQ2R[2]\ : NOR2
      port map(A => N_69, B => \DelayCnt_i[2]\, Y => N_72);
    
    \CycCnt_RNO_0[6]\ : AOI1
      port map(A => N_47, B => \CycCnt[5]_net_1\, C => 
        \CycCnt[6]_net_1\, Y => N_192);
    
    \CycCnt[9]\ : DFN1E1C0
      port map(D => CycCnt_n9, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[9]_net_1\);
    
    \Phase2Cnt_RNIKGGK[2]\ : OR3B
      port map(A => \Phase2Cnt[0]_net_1\, B => 
        \Phase2Cnt[2]_net_1\, C => \Phase2Cnt[1]_net_1\, Y => 
        N_73);
    
    \CycCnt_RNO[7]\ : XA1C
      port map(A => \CycCnt[7]_net_1\, B => N_68, C => 
        \PrState[4]_net_1\, Y => N_25_i_0);
    
    \PrState_RNO_0[0]\ : OR3A
      port map(A => \PrState_ns_0_0_a2_0_0[4]\, B => 
        \CycCnt[9]_net_1\, C => N_74, Y => N_92);
    
    \Phase2Cnt_RNO[2]\ : NOR3A
      port map(A => \PrState[1]_net_1\, B => N_116, C => N_117, Y
         => N_33);
    
    \DelayCnt_RNIRTH[1]\ : OR2B
      port map(A => \DelayCnt[1]_net_1\, B => \DelayCnt[0]_net_1\, 
        Y => N_69);
    
    \PrState_RNO_4[2]\ : NOR3A
      port map(A => lvdsFifoRowRdOut, B => \DelayCnt[0]_net_1\, C
         => \DelayCnt[1]_net_1\, Y => \PrState_ns_0_0_a2_0_2[2]\);
    
    \DelayCnt_RNO[1]\ : XA1
      port map(A => \DelayCnt[0]_net_1\, B => \DelayCnt[1]_net_1\, 
        C => \PrState[3]_net_1\, Y => N_35);
    
    \DelayCnt_RNI0II[4]\ : OR2B
      port map(A => \DelayCnt_i[2]\, B => \DelayCnt[4]_net_1\, Y
         => \PrState_ns_0_i_a2_0[1]\);
    
    \Phase2Cnt_RNO[1]\ : XA1
      port map(A => \Phase2Cnt[0]_net_1\, B => 
        \Phase2Cnt[1]_net_1\, C => \PrState[1]_net_1\, Y => N_31);
    
    \CycCnt[8]\ : DFN1E1C0
      port map(D => N_27_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[8]_net_1\);
    
    \CycCnt[5]\ : DFN1E1C0
      port map(D => N_21, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[5]_net_1\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \CycCnt_RNO[4]\ : XA1B
      port map(A => \CycCnt[4]_net_1\, B => N_46, C => 
        \PrState[4]_net_1\, Y => N_19);
    
    \CycCnt[0]\ : DFN1E1C0
      port map(D => CycCnt_n0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[0]_net_1\);
    
    \PrState_RNO_1[3]\ : OR3
      port map(A => \DelayCnt[0]_net_1\, B => \DelayCnt[1]_net_1\, 
        C => \PrState[4]_net_1\, Y => \PrState_ns_0_i_a2_1[1]\);
    
    \PrState_RNILTDS[1]\ : OR2A
      port map(A => \PrState[1]_net_1\, B => N_73, Y => N_78);
    
    \CycCnt_RNO[9]\ : XA1C
      port map(A => \CycCnt[9]_net_1\, B => N_74, C => 
        \PrState[4]_net_1\, Y => CycCnt_n9);
    
    \PrState[1]\ : DFN1C0
      port map(D => \PrState_ns[3]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \PrState[1]_net_1\);
    
    \DelayCnt_RNO[4]\ : NOR2A
      port map(A => \PrState[3]_net_1\, B => N_79_i, Y => N_41);
    
    \CycCnt_RNIUQ251[6]\ : OR3C
      port map(A => \CycCnt[5]_net_1\, B => N_47, C => 
        \CycCnt[6]_net_1\, Y => N_68);
    
    \CycCnt_RNO[6]\ : NOR3A
      port map(A => N_68, B => N_192, C => \PrState[4]_net_1\, Y
         => N_23);
    
    \PrState_RNO_0[2]\ : AOI1B
      port map(A => N_78, B => N_67, C => lvdsFifoRowRdOut, Y => 
        \PrState_ns_0_0_a2_0[2]\);
    
    \PrState_RNI7QQF[3]\ : NOR2
      port map(A => \PrState[4]_net_1\, B => \PrState[3]_net_1\, 
        Y => N_150);
    
    \CycCnt[2]\ : DFN1E1C0
      port map(D => N_15, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[2]_net_1\);
    
    \CycCnt_RNO[3]\ : XA1B
      port map(A => \CycCnt[3]_net_1\, B => N_177, C => 
        \PrState[4]_net_1\, Y => N_17);
    
    \CycCnt_RNO[2]\ : XA1B
      port map(A => \CycCnt[2]_net_1\, B => N_44, C => 
        \PrState[4]_net_1\, Y => N_15);
    
    \PrState_RNO[2]\ : AO1B
      port map(A => \PrState_ns_0_0_a2_0[2]\, B => N_129, C => 
        N_186_i, Y => \PrState_ns[2]\);
    
    \PrState_RNI57ON[0]\ : NOR3
      port map(A => \PrState[0]_net_1\, B => \PrState[2]_net_1\, 
        C => \PrState[3]_net_1\, Y => CycCntlde_0_a2_0_0);
    
    \CycCnt_RNO[0]\ : NOR2
      port map(A => \PrState[4]_net_1\, B => \CycCnt[0]_net_1\, Y
         => CycCnt_n0);
    
    \DelayCnt[2]\ : DFN1P0
      port map(D => N_37, CLK => PLL_Test1_0_Sys_66M_Clk, PRE => 
        PLL_Test1_0_SysRst_O, Q => \DelayCnt_i[2]\);
    
    \PrState_RNO_2[3]\ : OR2A
      port map(A => lvdsFifoRowRdOut, B => N_150, Y => 
        \PrState_ns_0_i_0[1]\);
    
    \CycCnt[6]\ : DFN1E1C0
      port map(D => N_23, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[6]_net_1\);
    
    \PrState_RNO_0[1]\ : NOR2B
      port map(A => \PrState[1]_net_1\, B => lvdsFifoRowRdOut, Y
         => \PrState_ns_0_0_a2_0[3]\);
    
    \Phase2Cnt[2]\ : DFN1C0
      port map(D => N_33, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase2Cnt[2]_net_1\);
    
    \Phase1Cnt[0]\ : DFN1C0
      port map(D => NxState_0_sqmuxa, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \Phase1Cnt[0]_net_1\);
    
    \DelayCnt[1]\ : DFN1C0
      port map(D => N_35, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \DelayCnt[1]_net_1\);
    
    \PrState_RNO_0[3]\ : OR2
      port map(A => \DelayCnt[3]_net_1\, B => 
        \PrState_ns_0_i_a2_0[1]\, Y => \PrState_ns_0_i_a2_0_0[1]\);
    
    \CycCnt[3]\ : DFN1E1C0
      port map(D => N_17, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[3]_net_1\);
    
    \Phase2Cnt_RNO[0]\ : NOR2A
      port map(A => \PrState[1]_net_1\, B => \Phase2Cnt[0]_net_1\, 
        Y => Phase2Cnt_n0);
    
    \DelayCnt[3]\ : DFN1C0
      port map(D => N_39, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \DelayCnt[3]_net_1\);
    
    \PrState_RNO[1]\ : AO1B
      port map(A => \PrState_ns_0_0_a2_0[3]\, B => N_73, C => 
        N_90, Y => \PrState_ns[3]\);
    
    \PrState[4]\ : DFN1P0
      port map(D => \PrState_RNO_3[4]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, PRE => PLL_Test1_0_SysRst_O, Q
         => \PrState[4]_net_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \CycCnt_RNO[1]\ : XA1B
      port map(A => \CycCnt[0]_net_1\, B => \CycCnt[1]_net_1\, C
         => \PrState[4]_net_1\, Y => N_13);
    
    \CycCnt[1]\ : DFN1E1C0
      port map(D => N_13, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[1]_net_1\);
    
    \Phase1Cnt_RNI2JME[0]\ : OR2B
      port map(A => \PrState[2]_net_1\, B => \Phase1Cnt[0]_net_1\, 
        Y => N_67);
    
    \DelayCnt_RNO[2]\ : XAI1
      port map(A => \DelayCnt_i[2]\, B => N_69, C => 
        \PrState[3]_net_1\, Y => N_37);
    
    \DelayCnt[4]\ : DFN1C0
      port map(D => N_41, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \DelayCnt[4]_net_1\);
    
    \DelayCnt_RNO[3]\ : XA1
      port map(A => \DelayCnt[3]_net_1\, B => N_72, C => 
        \PrState[3]_net_1\, Y => N_39);
    
    \Phase2Cnt[1]\ : DFN1C0
      port map(D => N_31, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase2Cnt[1]_net_1\);
    
    \DelayCnt[0]\ : DFN1C0
      port map(D => DelayCnt_n0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \DelayCnt[0]_net_1\);
    
    \CycCnt_RNIKSCA1[7]\ : OR2A
      port map(A => \CycCnt[7]_net_1\, B => N_68, Y => N_70);
    
    \PrState[0]\ : DFN1C0
      port map(D => \PrState_ns[4]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \PrState[0]_net_1\);
    
    \Phase1Cnt_RNI2JME_0[0]\ : NOR2A
      port map(A => \PrState[2]_net_1\, B => \Phase1Cnt[0]_net_1\, 
        Y => NxState_0_sqmuxa);
    
    \CycCnt_RNIVEIA[1]\ : NOR2B
      port map(A => \CycCnt[1]_net_1\, B => \CycCnt[0]_net_1\, Y
         => N_44);
    
    \CycCnt[4]\ : DFN1E1C0
      port map(D => N_19, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[4]_net_1\);
    
    \PrState_RNO[3]\ : OA1B
      port map(A => \PrState_ns_0_i_a2_0_0[1]\, B => 
        \PrState_ns_0_i_a2_1[1]\, C => \PrState_ns_0_i_0[1]\, Y
         => N_7);
    
    \Phase2Cnt_RNO_0[2]\ : AOI1
      port map(A => \Phase2Cnt[1]_net_1\, B => 
        \Phase2Cnt[0]_net_1\, C => \Phase2Cnt[2]_net_1\, Y => 
        N_116);
    
    \CycCnt[7]\ : DFN1E1C0
      port map(D => N_25_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[7]_net_1\);
    
    \PrState[3]\ : DFN1C0
      port map(D => N_7, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \PrState[3]_net_1\);
    
    \CycCnt_RNIGSRF[2]\ : NOR2B
      port map(A => N_44, B => \CycCnt[2]_net_1\, Y => N_177);
    
    \CycCnt_RNIB2NF1[8]\ : OR2A
      port map(A => \CycCnt[8]_net_1\, B => N_70, Y => N_74);
    
    \PrState_RNO_1[2]\ : OR3A
      port map(A => N_67, B => \CycCnt[9]_net_1\, C => N_74, Y
         => N_129);
    
    \PrState_RNO[0]\ : AO1B
      port map(A => \PrState[0]_net_1\, B => lvdsFifoRowRdOut, C
         => N_92, Y => \PrState_ns[4]\);
    
    \Phase2Cnt_RNO_1[2]\ : NOR3C
      port map(A => \Phase2Cnt[0]_net_1\, B => 
        \Phase2Cnt[2]_net_1\, C => \Phase2Cnt[1]_net_1\, Y => 
        N_117);
    
    \PrState_RNO_0[4]\ : NOR3
      port map(A => \PrState[0]_net_1\, B => \PrState[2]_net_1\, 
        C => \PrState[1]_net_1\, Y => \PrState_ns_i_0_a2_0[0]\);
    
    \PrState_RNIT46K1[4]\ : AO1A
      port map(A => N_73, B => CycCntlde_0_a2_0_0, C => 
        \PrState[4]_net_1\, Y => CycCnte);
    
    \CycCnt_RNIL3FQ[4]\ : NOR2B
      port map(A => N_46, B => \CycCnt[4]_net_1\, Y => N_47);
    
    \CycCnt_RNO[5]\ : XA1B
      port map(A => \CycCnt[5]_net_1\, B => N_47, C => 
        \PrState[4]_net_1\, Y => N_21);
    
    \CycCnt_RNO[8]\ : XA1C
      port map(A => \CycCnt[8]_net_1\, B => N_70, C => 
        \PrState[4]_net_1\, Y => N_27_i_0);
    
    \PrState_RNO_2[2]\ : OR3B
      port map(A => \PrState_ns_0_0_a2_0_0[2]\, B => 
        \PrState_ns_0_0_a2_0_2[2]\, C => \PrState_ns_0_i_a2_0[1]\, 
        Y => N_186_i);
    
    \PrState_RNO_1[1]\ : OR2B
      port map(A => NxState_0_sqmuxa, B => lvdsFifoRowRdOut, Y
         => N_90);
    
    \Phase2Cnt[0]\ : DFN1C0
      port map(D => Phase2Cnt_n0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \Phase2Cnt[0]_net_1\);
    
    \PrState_RNO[4]\ : AOI1
      port map(A => \PrState_ns_i_0_a2_0[0]\, B => N_150, C => 
        lvdsFifoRowRdOut, Y => \PrState_RNO_3[4]\);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    \PrState_RNO_1[0]\ : NOR2A
      port map(A => lvdsFifoRowRdOut, B => N_78, Y => 
        \PrState_ns_0_0_a2_0_0[4]\);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    \DelayCnt_RNO[0]\ : NOR2A
      port map(A => \PrState[3]_net_1\, B => \DelayCnt[0]_net_1\, 
        Y => DelayCnt_n0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3;
use proasic3.all;

entity WaveGenSingleZ15 is

    port( Main_ctl4SD_0_Fifo_wr   : out   std_logic;
          PLL_Test1_0_SysRst_O    : in    std_logic;
          PLL_Test1_0_Sys_66M_Clk : in    std_logic;
          FifoRowRdOut_1          : in    std_logic;
          FifoRowRdOut_0          : in    std_logic
        );

end WaveGenSingleZ15;

architecture DEF_ARCH of WaveGenSingleZ15 is 

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component XA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component XA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OAI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component XA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XAI1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \PrState_ns_0_i_0[3]\, \Phase1Cnt_RNIIFV7[0]_net_1\, 
        \PrState[1]_net_1\, \PrState_ns_0_i_0[1]\, N_181, 
        \PrState_ns_i_0_a3_1[0]\, \PrState[0]_net_1\, 
        \PrState[2]_net_1\, \PrState_ns_0_i_a3_0_0[1]\, 
        \DelayCnt_i_0[3]\, \DelayCnt[2]_net_1\, 
        \PrState[4]_net_1\, \PrState_ns_0_0_a3_1_2_0[2]\, 
        \PrState[3]_net_1\, CycCntlde_0_a3_1, N_33, 
        \DelayCnt[0]_net_1\, \DelayCnt[1]_net_1\, N_35, N_163, 
        N_17, N_180, N_14, N_29_i_0, \CycCnt[8]_net_1\, N_45, 
        N_27_i_0, \CycCnt[7]_net_1\, N_43, N_25, N_175, N_23, 
        \CycCnt[5]_net_1\, N_161, N_21, \CycCnt[0]_net_1\, 
        \CycCnt[1]_net_1\, \PrState_ns_0_0_a3_0[2]\, N_68, 
        \CycCnt[9]_net_1\, N_162, N_172, \PrState_ns_0_0_0_tz[2]\, 
        \PrState_ns_0_0_a3_0_0[2]\, \Phase1Cnt[0]_net_1\, 
        \PrState_ns[2]\, DelayCnt_n0, \Phase2Cnt[1]_net_1\, 
        N_159_i_0, N_5, N_7, \PrState_RNO_0[4]_net_1\, 
        \PrState_ns[4]\, N_37, N_166, N_13, N_12, 
        \CycCnt[3]_net_1\, N_38, \CycCnt[2]_net_1\, N_9, 
        \CycCnt[4]_net_1\, N_183, N_182, \CycCnt[6]_net_1\, 
        CycCnt_n9, CycCnte, CycCnt_n0, \GND\, \VCC\, GND_0, VCC_0
         : std_logic;

begin 


    WFO : DFN1C0
      port map(D => \PrState[2]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => Main_ctl4SD_0_Fifo_wr);
    
    \PrState_RNITT97[0]\ : NOR3
      port map(A => \PrState[2]_net_1\, B => \PrState[0]_net_1\, 
        C => \PrState[3]_net_1\, Y => CycCntlde_0_a3_1);
    
    \PrState[2]\ : DFN1C0
      port map(D => \PrState_ns[2]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \PrState[2]_net_1\);
    
    \PrState_RNO_3[2]\ : OR2B
      port map(A => \PrState[2]_net_1\, B => \Phase1Cnt[0]_net_1\, 
        Y => \PrState_ns_0_0_a3_0_0[2]\);
    
    \Phase1Cnt_RNIIFV7[0]\ : NOR2A
      port map(A => \PrState[2]_net_1\, B => \Phase1Cnt[0]_net_1\, 
        Y => \Phase1Cnt_RNIIFV7[0]_net_1\);
    
    \CycCnt_RNO_0[6]\ : AOI1
      port map(A => N_161, B => \CycCnt[5]_net_1\, C => 
        \CycCnt[6]_net_1\, Y => N_175);
    
    \CycCnt[9]\ : DFN1E1C0
      port map(D => CycCnt_n9, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[9]_net_1\);
    
    \CycCnt_RNO[7]\ : XA1C
      port map(A => \CycCnt[7]_net_1\, B => N_43, C => 
        \PrState[4]_net_1\, Y => N_27_i_0);
    
    \PrState_RNO_0[0]\ : OR3A
      port map(A => \PrState_ns_0_0_a3_0[2]\, B => 
        \CycCnt[9]_net_1\, C => N_162, Y => N_172);
    
    \DelayCnt_RNO_0[3]\ : NOR2A
      port map(A => \DelayCnt[2]_net_1\, B => N_163, Y => N_166);
    
    \CycCnt_RNI2NI3[3]\ : NOR2B
      port map(A => N_12, B => \CycCnt[3]_net_1\, Y => N_13);
    
    \DelayCnt_RNO[1]\ : XA1
      port map(A => \DelayCnt[0]_net_1\, B => \DelayCnt[1]_net_1\, 
        C => \PrState[3]_net_1\, Y => N_33);
    
    \PrState_RNIIBDH[1]\ : NOR3B
      port map(A => \PrState[1]_net_1\, B => FifoRowRdOut_0, C
         => N_180, Y => \PrState_ns_0_0_a3_0[2]\);
    
    \Phase2Cnt_RNO[1]\ : XA1
      port map(A => N_159_i_0, B => \Phase2Cnt[1]_net_1\, C => 
        \PrState[1]_net_1\, Y => N_7);
    
    \CycCnt[8]\ : DFN1E1C0
      port map(D => N_29_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[8]_net_1\);
    
    \CycCnt[5]\ : DFN1E1C0
      port map(D => N_23, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[5]_net_1\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \CycCnt_RNO[4]\ : XA1B
      port map(A => \CycCnt[4]_net_1\, B => N_13, C => 
        \PrState[4]_net_1\, Y => N_9);
    
    \CycCnt[0]\ : DFN1E1C0
      port map(D => CycCnt_n0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[0]_net_1\);
    
    \PrState_RNO_1[3]\ : NOR2B
      port map(A => FifoRowRdOut_0, B => N_181, Y => 
        \PrState_ns_0_i_0[1]\);
    
    \PrState_RNIG7UK[4]\ : AO1A
      port map(A => N_180, B => CycCntlde_0_a3_1, C => 
        \PrState[4]_net_1\, Y => CycCnte);
    
    \CycCnt_RNO[9]\ : XA1C
      port map(A => \CycCnt[9]_net_1\, B => N_162, C => 
        \PrState[4]_net_1\, Y => CycCnt_n9);
    
    \PrState[1]\ : DFN1C0
      port map(D => N_17, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \PrState[1]_net_1\);
    
    \CycCnt_RNO[6]\ : NOR3A
      port map(A => N_43, B => N_175, C => \PrState[4]_net_1\, Y
         => N_25);
    
    \DelayCnt_RNIB2J4[1]\ : OR2B
      port map(A => \DelayCnt[1]_net_1\, B => \DelayCnt[0]_net_1\, 
        Y => N_163);
    
    \PrState_RNO_0[2]\ : OA1A
      port map(A => \PrState_ns_0_0_a3_1_2_0[2]\, B => N_163, C
         => \PrState_ns_0_0_a3_0_0[2]\, Y => 
        \PrState_ns_0_0_0_tz[2]\);
    
    \CycCnt_RNIKE77[7]\ : OR2A
      port map(A => \CycCnt[7]_net_1\, B => N_43, Y => N_45);
    
    \CycCnt[2]\ : DFN1E1C0
      port map(D => N_182, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[2]_net_1\);
    
    \CycCnt_RNO[3]\ : XA1B
      port map(A => \CycCnt[3]_net_1\, B => N_12, C => 
        \PrState[4]_net_1\, Y => N_183);
    
    \CycCnt_RNO[2]\ : XA1B
      port map(A => \CycCnt[2]_net_1\, B => N_38, C => 
        \PrState[4]_net_1\, Y => N_182);
    
    \CycCnt_RNIM2A6[6]\ : OR3C
      port map(A => \CycCnt[5]_net_1\, B => N_161, C => 
        \CycCnt[6]_net_1\, Y => N_43);
    
    \PrState_RNO[2]\ : AO1C
      port map(A => \PrState_ns_0_0_0_tz[2]\, B => FifoRowRdOut_1, 
        C => N_68, Y => \PrState_ns[2]\);
    
    \CycCnt_RNO[0]\ : NOR2
      port map(A => \PrState[4]_net_1\, B => \CycCnt[0]_net_1\, Y
         => CycCnt_n0);
    
    \DelayCnt[2]\ : DFN1C0
      port map(D => N_35, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \DelayCnt[2]_net_1\);
    
    \CycCnt[6]\ : DFN1E1C0
      port map(D => N_25, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[6]_net_1\);
    
    \PrState_RNO_0[1]\ : OAI1
      port map(A => \Phase1Cnt_RNIIFV7[0]_net_1\, B => 
        \PrState[1]_net_1\, C => FifoRowRdOut_0, Y => 
        \PrState_ns_0_i_0[3]\);
    
    \Phase1Cnt[0]\ : DFN1C0
      port map(D => \Phase1Cnt_RNIIFV7[0]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \Phase1Cnt[0]_net_1\);
    
    \DelayCnt[1]\ : DFN1C0
      port map(D => N_33, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \DelayCnt[1]_net_1\);
    
    \CycCnt_RNITMF4[4]\ : NOR2B
      port map(A => N_13, B => \CycCnt[4]_net_1\, Y => N_161);
    
    \PrState_RNO_0[3]\ : NOR3
      port map(A => \DelayCnt_i_0[3]\, B => \DelayCnt[2]_net_1\, 
        C => \PrState[4]_net_1\, Y => \PrState_ns_0_i_a3_0_0[1]\);
    
    \CycCnt[3]\ : DFN1E1C0
      port map(D => N_183, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[3]_net_1\);
    
    \Phase2Cnt_RNO[0]\ : NOR2A
      port map(A => \PrState[1]_net_1\, B => N_159_i_0, Y => N_5);
    
    \DelayCnt[3]\ : DFN1P0
      port map(D => N_37, CLK => PLL_Test1_0_Sys_66M_Clk, PRE => 
        PLL_Test1_0_SysRst_O, Q => \DelayCnt_i_0[3]\);
    
    \CycCnt_RNIJU48[8]\ : OR2A
      port map(A => \CycCnt[8]_net_1\, B => N_45, Y => N_162);
    
    \PrState_RNO[1]\ : OA1B
      port map(A => \Phase1Cnt_RNIIFV7[0]_net_1\, B => N_180, C
         => \PrState_ns_0_i_0[3]\, Y => N_17);
    
    \PrState[4]\ : DFN1P0
      port map(D => \PrState_RNO_0[4]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, PRE => PLL_Test1_0_SysRst_O, Q
         => \PrState[4]_net_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \CycCnt_RNO[1]\ : XA1B
      port map(A => \CycCnt[0]_net_1\, B => \CycCnt[1]_net_1\, C
         => \PrState[4]_net_1\, Y => N_21);
    
    \CycCnt[1]\ : DFN1E1C0
      port map(D => N_21, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[1]_net_1\);
    
    \CycCnt_RNIF3P1[1]\ : NOR2B
      port map(A => \CycCnt[1]_net_1\, B => \CycCnt[0]_net_1\, Y
         => N_38);
    
    \DelayCnt_RNO[2]\ : XA1A
      port map(A => \DelayCnt[2]_net_1\, B => N_163, C => 
        \PrState[3]_net_1\, Y => N_35);
    
    \Phase2Cnt_RNI7A6B[1]\ : OR2A
      port map(A => \Phase2Cnt[1]_net_1\, B => N_159_i_0, Y => 
        N_180);
    
    \DelayCnt_RNO[3]\ : XAI1A
      port map(A => \DelayCnt_i_0[3]\, B => N_166, C => 
        \PrState[3]_net_1\, Y => N_37);
    
    \Phase2Cnt[1]\ : DFN1C0
      port map(D => N_7, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase2Cnt[1]_net_1\);
    
    \DelayCnt[0]\ : DFN1C0
      port map(D => DelayCnt_n0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \DelayCnt[0]_net_1\);
    
    \PrState[0]\ : DFN1C0
      port map(D => \PrState_ns[4]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \PrState[0]_net_1\);
    
    \PrState_RNINUR4[3]\ : OR2
      port map(A => \PrState[4]_net_1\, B => \PrState[3]_net_1\, 
        Y => N_181);
    
    \CycCnt_RNI8RL2[2]\ : NOR2B
      port map(A => N_38, B => \CycCnt[2]_net_1\, Y => N_12);
    
    \CycCnt[4]\ : DFN1E1C0
      port map(D => N_9, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[4]_net_1\);
    
    \PrState_RNO[3]\ : OA1A
      port map(A => \PrState_ns_0_i_a3_0_0[1]\, B => N_163, C => 
        \PrState_ns_0_i_0[1]\, Y => N_14);
    
    \CycCnt[7]\ : DFN1E1C0
      port map(D => N_27_i_0, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[7]_net_1\);
    
    \PrState[3]\ : DFN1C0
      port map(D => N_14, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \PrState[3]_net_1\);
    
    \PrState_RNO_1[2]\ : OAI1
      port map(A => \CycCnt[9]_net_1\, B => N_162, C => 
        \PrState_ns_0_0_a3_0[2]\, Y => N_68);
    
    \PrState_RNO[0]\ : AO1B
      port map(A => \PrState[0]_net_1\, B => FifoRowRdOut_1, C
         => N_172, Y => \PrState_ns[4]\);
    
    \PrState_RNO_0[4]\ : OR3
      port map(A => \PrState[1]_net_1\, B => \PrState[0]_net_1\, 
        C => \PrState[2]_net_1\, Y => \PrState_ns_i_0_a3_1[0]\);
    
    \CycCnt_RNO[5]\ : XA1B
      port map(A => \CycCnt[5]_net_1\, B => N_161, C => 
        \PrState[4]_net_1\, Y => N_23);
    
    \CycCnt_RNO[8]\ : XA1C
      port map(A => \CycCnt[8]_net_1\, B => N_45, C => 
        \PrState[4]_net_1\, Y => N_29_i_0);
    
    \PrState_RNO_2[2]\ : NOR3A
      port map(A => \PrState[3]_net_1\, B => \DelayCnt_i_0[3]\, C
         => \DelayCnt[2]_net_1\, Y => 
        \PrState_ns_0_0_a3_1_2_0[2]\);
    
    \Phase2Cnt[0]\ : DFN1C0
      port map(D => N_5, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => N_159_i_0);
    
    \PrState_RNO[4]\ : OA1B
      port map(A => N_181, B => \PrState_ns_i_0_a3_1[0]\, C => 
        FifoRowRdOut_1, Y => \PrState_RNO_0[4]_net_1\);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    \DelayCnt_RNO[0]\ : NOR2A
      port map(A => \PrState[3]_net_1\, B => \DelayCnt[0]_net_1\, 
        Y => DelayCnt_n0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3;
use proasic3.all;

entity WaveGenSingleZ13 is

    port( PLL_Test1_0_SysRst_O    : in    std_logic;
          PLL_Test1_0_Sys_66M_Clk : in    std_logic;
          FifoRowRdOut            : in    std_logic;
          Data2Fifo_0_sqmuxa      : out   std_logic;
          FifoRowRdOut_1          : in    std_logic;
          FifoRowRdOut_0          : in    std_logic;
          Data2Fifo_0_sqmuxa_0    : out   std_logic;
          CMOS_DrvX_0_SDramEn_0   : in    std_logic;
          Data2Fifo_0_sqmuxa_1    : out   std_logic
        );

end WaveGenSingleZ13;

architecture DEF_ARCH of WaveGenSingleZ13 is 

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component XA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1D
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component NOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal Data2fifoEN, \PrState_ns_i_0_a2_0[0]\, 
        \PrState[1]_net_1\, \PrState[2]_net_1\, 
        \PrState_ns_0_i_0[1]\, N_41, \PrState[3]_net_1\, 
        \PrState_ns_0_0_o2_6[2]\, \PrState_ns_0_0_o2_1[2]\, 
        \PrState_ns_0_0_o2_0[2]\, N_29, \PrState_ns_0_0_o2_5[2]\, 
        \CycCnt[4]_net_1\, \CycCnt[2]_net_1\, 
        \PrState_ns_0_0_o2_3[2]\, \CycCnt[6]_net_1\, 
        \CycCnt[8]_net_1\, \CycCnt[5]_net_1\, \CycCnt[7]_net_1\, 
        \CycCnt[3]_net_1\, \CycCnt[9]_net_1\, 
        \PrState_ns_0_i_a2_2[1]\, \DelayCnt[1]_net_1\, 
        \DelayCnt[3]_net_1\, \PrState_ns_0_i_a2_1[1]\, 
        \DelayCnt[0]_net_1\, \DelayCnt[2]_net_1\, 
        \PrState_ns_0_0_a2_1_2_1[2]\, CycCntlde_0_a2_1, 
        \PrState[0]_net_1\, N_175, N_173, N_17, N_19, N_26, N_177, 
        \CycCnt[0]_net_1\, \CycCnt[1]_net_1\, N_178, N_9, N_22, 
        N_179, N_193, N_24, N_13, N_15, N_197, N_183, N_180, 
        N_181, N_184, N_11, \PrState_ns_0_0_0_tz[2]\, DelayCnt_n0, 
        \PrState_ns_0_0_a2_0_0[2]\, \Phase1Cnt[0]_net_1\, 
        \PrState_ns[2]\, N_45, \Phase2Cnt[1]_net_1\, N_159_i_0, 
        N_5, N_7, N_14, N_27, N_39, N_21, N_28, CycCnt_n0, N_185, 
        N_43_2, CycCnt_n9, \PrState_ns[4]\, N_170, 
        \PrState_RNO_1[4]\, CycCnte, \GND\, \VCC\, GND_0, VCC_0
         : std_logic;

begin 


    WFO : DFN1C0
      port map(D => \PrState[2]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => Data2fifoEN);
    
    \PrState[2]\ : DFN1C0
      port map(D => \PrState_ns[2]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \PrState[2]_net_1\);
    
    \PrState_RNO_3[2]\ : OR2B
      port map(A => \PrState[2]_net_1\, B => \Phase1Cnt[0]_net_1\, 
        Y => \PrState_ns_0_0_a2_0_0[2]\);
    
    \CycCnt_RNIOKF7[7]\ : NOR2B
      port map(A => \CycCnt[5]_net_1\, B => \CycCnt[7]_net_1\, Y
         => \PrState_ns_0_0_o2_1[2]\);
    
    \CycCnt_RNO_0[6]\ : AO1A
      port map(A => N_24, B => \CycCnt[5]_net_1\, C => 
        \CycCnt[6]_net_1\, Y => N_197);
    
    \CycCnt[9]\ : DFN1E1C0
      port map(D => CycCnt_n9, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[9]_net_1\);
    
    WFO_RNI8L1B_0 : NOR2B
      port map(A => Data2fifoEN, B => CMOS_DrvX_0_SDramEn_0, Y
         => Data2Fifo_0_sqmuxa_0);
    
    \CycCnt_RNO_0[4]\ : AO1A
      port map(A => N_22, B => \CycCnt[3]_net_1\, C => 
        \CycCnt[4]_net_1\, Y => N_193);
    
    WFO_RNI8L1B : NOR2B
      port map(A => Data2fifoEN, B => CMOS_DrvX_0_SDramEn_0, Y
         => Data2Fifo_0_sqmuxa_1);
    
    \CycCnt_RNO[7]\ : XA1C
      port map(A => \CycCnt[7]_net_1\, B => N_183, C => N_41, Y
         => N_180);
    
    \PrState_RNO_0[0]\ : OR3C
      port map(A => \PrState_ns_0_0_o2_5[2]\, B => 
        \PrState_ns_0_0_o2_6[2]\, C => N_175, Y => N_170);
    
    \DelayCnt_RNO_0[3]\ : NOR2B
      port map(A => N_26, B => \DelayCnt[2]_net_1\, Y => N_28);
    
    \DelayCnt_RNO[1]\ : XA1
      port map(A => \DelayCnt[0]_net_1\, B => \DelayCnt[1]_net_1\, 
        C => \PrState[3]_net_1\, Y => N_17);
    
    \Phase2Cnt_RNO[1]\ : XA1
      port map(A => N_159_i_0, B => \Phase2Cnt[1]_net_1\, C => 
        \PrState[1]_net_1\, Y => N_7);
    
    \CycCnt_RNILI5B[2]\ : OR2A
      port map(A => \CycCnt[2]_net_1\, B => N_29, Y => N_22);
    
    \CycCnt[8]\ : DFN1E1C0
      port map(D => N_181, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[8]_net_1\);
    
    \CycCnt[5]\ : DFN1E1C0
      port map(D => N_13, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[5]_net_1\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \CycCnt_RNO[4]\ : NOR3B
      port map(A => N_193, B => N_24, C => N_41, Y => N_179);
    
    \CycCnt[0]\ : DFN1E1C0
      port map(D => CycCnt_n0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[0]_net_1\);
    
    \CycCnt_RNIOKF7[9]\ : NOR2A
      port map(A => \CycCnt[3]_net_1\, B => \CycCnt[9]_net_1\, Y
         => \PrState_ns_0_0_o2_0[2]\);
    
    \PrState_RNO_1[3]\ : NOR2
      port map(A => \DelayCnt[0]_net_1\, B => \DelayCnt[2]_net_1\, 
        Y => \PrState_ns_0_i_a2_1[1]\);
    
    \CycCnt_RNO[9]\ : XA1
      port map(A => \CycCnt[9]_net_1\, B => N_185, C => N_43_2, Y
         => CycCnt_n9);
    
    \PrState_RNIIMB2[4]\ : AO1D
      port map(A => CycCntlde_0_a2_1, B => N_173, C => N_41, Y
         => CycCnte);
    
    \PrState[1]\ : DFN1C0
      port map(D => N_14, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \PrState[1]_net_1\);
    
    \CycCnt_RNO_0[9]\ : NOR2B
      port map(A => N_184, B => \CycCnt[8]_net_1\, Y => N_185);
    
    \CycCnt_RNO[6]\ : NOR3B
      port map(A => N_197, B => N_183, C => N_41, Y => N_15);
    
    \DelayCnt_RNILOE6[0]\ : NOR2B
      port map(A => \DelayCnt[1]_net_1\, B => \DelayCnt[0]_net_1\, 
        Y => N_26);
    
    \CycCnt_RNI8JKI[4]\ : OR3B
      port map(A => \CycCnt[3]_net_1\, B => \CycCnt[4]_net_1\, C
         => N_22, Y => N_24);
    
    \PrState_RNO_0[2]\ : AOI1B
      port map(A => \PrState_ns_0_0_a2_1_2_1[2]\, B => 
        DelayCnt_n0, C => \PrState_ns_0_0_a2_0_0[2]\, Y => 
        \PrState_ns_0_0_0_tz[2]\);
    
    \CycCnt[2]\ : DFN1E1C0
      port map(D => N_178, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[2]_net_1\);
    
    \CycCnt_RNO[3]\ : XA1C
      port map(A => \CycCnt[3]_net_1\, B => N_22, C => N_41, Y
         => N_9);
    
    \CycCnt_RNO[2]\ : XA1C
      port map(A => \CycCnt[2]_net_1\, B => N_29, C => N_41, Y
         => N_178);
    
    \PrState_RNO[2]\ : AO1C
      port map(A => \PrState_ns_0_0_0_tz[2]\, B => FifoRowRdOut_0, 
        C => N_45, Y => \PrState_ns[2]\);
    
    \CycCnt_RNO[0]\ : NOR2
      port map(A => N_41, B => \CycCnt[0]_net_1\, Y => CycCnt_n0);
    
    \DelayCnt[2]\ : DFN1C0
      port map(D => N_19, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \DelayCnt[2]_net_1\);
    
    \PrState_RNO_2[3]\ : OA1
      port map(A => N_41, B => \PrState[3]_net_1\, C => 
        FifoRowRdOut_0, Y => \PrState_ns_0_i_0[1]\);
    
    \CycCnt[6]\ : DFN1E1C0
      port map(D => N_15, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[6]_net_1\);
    
    \PrState_RNO_0[1]\ : NOR2B
      port map(A => \PrState[1]_net_1\, B => N_173, Y => N_39);
    
    \Phase1Cnt[0]\ : DFN1C0
      port map(D => N_27, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase1Cnt[0]_net_1\);
    
    \DelayCnt_RNIQ0N3[0]\ : NOR2A
      port map(A => \PrState[3]_net_1\, B => \DelayCnt[0]_net_1\, 
        Y => DelayCnt_n0);
    
    \DelayCnt[1]\ : DFN1C0
      port map(D => N_17, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \DelayCnt[1]_net_1\);
    
    WFO_RNI8L1B_1 : NOR2B
      port map(A => Data2fifoEN, B => CMOS_DrvX_0_SDramEn_0, Y
         => Data2Fifo_0_sqmuxa);
    
    \PrState_RNO_0[3]\ : NOR3B
      port map(A => \DelayCnt[1]_net_1\, B => \DelayCnt[3]_net_1\, 
        C => N_41, Y => \PrState_ns_0_i_a2_2[1]\);
    
    \CycCnt[3]\ : DFN1E1C0
      port map(D => N_9, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[3]_net_1\);
    
    \Phase2Cnt_RNO[0]\ : NOR2A
      port map(A => \PrState[1]_net_1\, B => N_159_i_0, Y => N_5);
    
    \DelayCnt[3]\ : DFN1C0
      port map(D => N_21, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \DelayCnt[3]_net_1\);
    
    \PrState_RNO[1]\ : OA1
      port map(A => N_27, B => N_39, C => FifoRowRdOut_1, Y => 
        N_14);
    
    \PrState[4]\ : DFN1P0
      port map(D => \PrState_RNO_1[4]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, PRE => PLL_Test1_0_SysRst_O, Q
         => N_41);
    
    \CycCnt_RNID8E7[1]\ : OR2B
      port map(A => \CycCnt[1]_net_1\, B => \CycCnt[0]_net_1\, Y
         => N_29);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \PrState_RNIE3F1[0]\ : NOR3
      port map(A => N_41, B => \PrState[3]_net_1\, C => 
        \PrState[0]_net_1\, Y => N_43_2);
    
    \CycCnt_RNO[1]\ : XA1B
      port map(A => \CycCnt[0]_net_1\, B => \CycCnt[1]_net_1\, C
         => N_41, Y => N_177);
    
    \CycCnt[1]\ : DFN1E1C0
      port map(D => N_177, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[1]_net_1\);
    
    \DelayCnt_RNO[2]\ : XA1
      port map(A => \DelayCnt[2]_net_1\, B => N_26, C => 
        \PrState[3]_net_1\, Y => N_19);
    
    \DelayCnt_RNO[3]\ : XA1
      port map(A => \DelayCnt[3]_net_1\, B => N_28, C => 
        \PrState[3]_net_1\, Y => N_21);
    
    \Phase2Cnt[1]\ : DFN1C0
      port map(D => N_7, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \Phase2Cnt[1]_net_1\);
    
    \CycCnt_RNIV34Q[6]\ : OR3B
      port map(A => \CycCnt[5]_net_1\, B => \CycCnt[6]_net_1\, C
         => N_24, Y => N_183);
    
    \DelayCnt[0]\ : DFN1C0
      port map(D => DelayCnt_n0, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \DelayCnt[0]_net_1\);
    
    \PrState[0]\ : DFN1C0
      port map(D => \PrState_ns[4]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \PrState[0]_net_1\);
    
    \CycCnt_RNIQSF7[6]\ : NOR2B
      port map(A => \CycCnt[6]_net_1\, B => \CycCnt[8]_net_1\, Y
         => \PrState_ns_0_0_o2_3[2]\);
    
    \PrState_RNI5LL4[1]\ : NOR3B
      port map(A => \PrState[1]_net_1\, B => FifoRowRdOut_0, C
         => N_173, Y => N_175);
    
    \CycCnt_RNICPUE[2]\ : NOR3C
      port map(A => \CycCnt[4]_net_1\, B => \CycCnt[2]_net_1\, C
         => \PrState_ns_0_0_o2_3[2]\, Y => 
        \PrState_ns_0_0_o2_5[2]\);
    
    \PrState_RNIC3F1[0]\ : OR3
      port map(A => \PrState[0]_net_1\, B => \PrState[3]_net_1\, 
        C => \PrState[2]_net_1\, Y => CycCntlde_0_a2_1);
    
    \CycCnt[4]\ : DFN1E1C0
      port map(D => N_179, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[4]_net_1\);
    
    \PrState_RNO[3]\ : AOI1B
      port map(A => \PrState_ns_0_i_a2_2[1]\, B => 
        \PrState_ns_0_i_a2_1[1]\, C => \PrState_ns_0_i_0[1]\, Y
         => N_11);
    
    \CycCnt[7]\ : DFN1E1C0
      port map(D => N_180, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CycCnte, Q => 
        \CycCnt[7]_net_1\);
    
    \PrState[3]\ : DFN1C0
      port map(D => N_11, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => \PrState[3]_net_1\);
    
    \CycCnt_RNITHDM[7]\ : NOR3B
      port map(A => \PrState_ns_0_0_o2_1[2]\, B => 
        \PrState_ns_0_0_o2_0[2]\, C => N_29, Y => 
        \PrState_ns_0_0_o2_6[2]\);
    
    \PrState_RNO_1[2]\ : AO1B
      port map(A => \PrState_ns_0_0_o2_6[2]\, B => 
        \PrState_ns_0_0_o2_5[2]\, C => N_175, Y => N_45);
    
    \PrState_RNO[0]\ : AO1B
      port map(A => FifoRowRdOut, B => \PrState[0]_net_1\, C => 
        N_170, Y => \PrState_ns[4]\);
    
    \PrState_RNO_0[4]\ : OR2
      port map(A => \PrState[1]_net_1\, B => \PrState[2]_net_1\, 
        Y => \PrState_ns_i_0_a2_0[0]\);
    
    \CycCnt_RNO[5]\ : XA1C
      port map(A => \CycCnt[5]_net_1\, B => N_24, C => N_41, Y
         => N_13);
    
    \CycCnt_RNIC2ST[7]\ : NOR2A
      port map(A => \CycCnt[7]_net_1\, B => N_183, Y => N_184);
    
    \Phase1Cnt_RNIUFK[0]\ : NOR2A
      port map(A => \PrState[2]_net_1\, B => \Phase1Cnt[0]_net_1\, 
        Y => N_27);
    
    \CycCnt_RNO[8]\ : XA1B
      port map(A => \CycCnt[8]_net_1\, B => N_184, C => N_41, Y
         => N_181);
    
    \PrState_RNO_2[2]\ : NOR3B
      port map(A => \DelayCnt[1]_net_1\, B => \DelayCnt[3]_net_1\, 
        C => \DelayCnt[2]_net_1\, Y => 
        \PrState_ns_0_0_a2_1_2_1[2]\);
    
    \Phase2Cnt[0]\ : DFN1C0
      port map(D => N_5, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, Q => N_159_i_0);
    
    \PrState_RNO[4]\ : OA1C
      port map(A => N_43_2, B => \PrState_ns_i_0_a2_0[0]\, C => 
        FifoRowRdOut, Y => \PrState_RNO_1[4]\);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    \Phase2Cnt_RNILSC[1]\ : OR2A
      port map(A => \Phase2Cnt[1]_net_1\, B => N_159_i_0, Y => 
        N_173);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3;
use proasic3.all;

entity Main_ctl4SD is

    port( intData2acc_RNIPB46                 : out   std_logic_vector(71 to 71);
          intData2acc_RNIFHV6                 : out   std_logic_vector(4 to 4);
          intData2acc_RNIEDV6                 : out   std_logic_vector(3 to 3);
          intData2acc_RNIITV6                 : out   std_logic_vector(7 to 7);
          intData2acc_RNIHPV6                 : out   std_logic_vector(6 to 6);
          intData2acc_RNIGLV6                 : out   std_logic_vector(5 to 5);
          intData2acc_RNI6J36                 : out   std_logic_vector(10 to 10);
          intData2acc_RNIK507                 : out   std_logic_vector(9 to 9);
          intData2acc_RNIJ107                 : out   std_logic_vector(8 to 8);
          intData2acc_RNI9J36                 : out   std_logic_vector(13 to 13);
          intData2acc_RNI8J36                 : out   std_logic_vector(12 to 12);
          intData2acc_RNI7J36                 : out   std_logic_vector(11 to 11);
          intData2acc_RNICJ36                 : out   std_logic_vector(16 to 16);
          intData2acc_RNIBJ36                 : out   std_logic_vector(15 to 15);
          intData2acc_RNIAJ36                 : out   std_logic_vector(14 to 14);
          intData2acc_RNIDJ36                 : out   std_logic_vector(17 to 17);
          intData2acc_RNIBN36                 : out   std_logic_vector(22 to 22);
          intData2acc_RNIAN36                 : out   std_logic_vector(21 to 21);
          intData2acc_RNIEN36                 : out   std_logic_vector(25 to 25);
          intData2acc_RNIDN36                 : out   std_logic_vector(24 to 24);
          intData2acc_RNITJS7                 : out   std_logic_vector(23 to 23);
          intData2acc_RNI2KS7                 : out   std_logic_vector(28 to 28);
          intData2acc_RNI1KS7                 : out   std_logic_vector(27 to 27);
          intData2acc_RNI0KS7                 : out   std_logic_vector(26 to 26);
          intData2acc_RNI4JV9                 : out   std_logic_vector(31 to 31);
          intData2acc_RNI3JV9                 : out   std_logic_vector(30 to 30);
          intData2acc_RNI9FV9                 : out   std_logic_vector(29 to 29);
          intData2acc_RNI5JV9                 : out   std_logic_vector(32 to 32);
          intData2acc_RNI8JV9                 : out   std_logic_vector(35 to 35);
          intData2acc_RNI6NV9                 : out   std_logic_vector(40 to 40);
          intData2acc_RNICJV9                 : out   std_logic_vector(39 to 39);
          intData2acc_RNIBJV9                 : out   std_logic_vector(38 to 38);
          intData2acc_RNI9NV9                 : out   std_logic_vector(43 to 43);
          intData2acc_RNI8NV9                 : out   std_logic_vector(42 to 42);
          intData2acc_RNI7NV9                 : out   std_logic_vector(41 to 41);
          intData2acc_RNICNV9                 : out   std_logic_vector(46 to 46);
          intData2acc_RNIBNV9                 : out   std_logic_vector(45 to 45);
          intData2acc_RNIANV9                 : out   std_logic_vector(44 to 44);
          intData2acc_RNIFNV9                 : out   std_logic_vector(49 to 49);
          intData2acc_RNIENV9                 : out   std_logic_vector(48 to 48);
          intData2acc_RNIDNV9                 : out   std_logic_vector(47 to 47);
          intData2acc_RNI9RV9                 : out   std_logic_vector(51 to 51);
          intData2acc_RNI8RV9                 : out   std_logic_vector(50 to 50);
          intData2acc_RNIERV9                 : out   std_logic_vector(57 to 57);
          intData2acc_RNIDRV9                 : out   std_logic_vector(56 to 56);
          intData2acc_RNIBVV9                 : out   std_logic_vector(61 to 61);
          intData2acc_RNIAVV9                 : out   std_logic_vector(60 to 60);
          intData2acc_RNIGRV9                 : out   std_logic_vector(59 downto 58);
          intData2acc_RNIEVV9                 : out   std_logic_vector(64 to 64);
          intData2acc_RNIDVV9                 : out   std_logic_vector(63 to 63);
          intData2acc_RNICVV9                 : out   std_logic_vector(62 to 62);
          intData2acc_RNIHVV9                 : out   std_logic_vector(67 to 67);
          intData2acc_RNIGVV9                 : out   std_logic_vector(66 to 66);
          intData2acc_RNIFVV9                 : out   std_logic_vector(65 to 65);
          intData2acc_RNID30A                 : out   std_logic_vector(70 to 70);
          intData2acc_RNIVOQA                 : out   std_logic_vector(0 to 0);
          intData2acc_RNI2BV9                 : out   std_logic_vector(18 to 18);
          intData2acc_RNI6JV9_0               : out   std_logic;
          intData2acc_RNI6JV9_3               : out   std_logic;
          intData2acc_RNI0TQA                 : out   std_logic_vector(1 to 1);
          intData2acc_RNI3BV9                 : out   std_logic_vector(19 to 19);
          intData2acc_RNI7JV9_0               : out   std_logic;
          intData2acc_RNI7JV9_3               : out   std_logic;
          intData2acc_RNI11RA                 : out   std_logic_vector(2 to 2);
          intData2acc_RNITEV9                 : out   std_logic_vector(20 to 20);
          pr_state_ns                         : in    std_logic_vector(8 to 8);
          intData2acc_RNIARV9                 : out   std_logic_vector(54 to 54);
          intData2acc_RNIBRV9_0               : out   std_logic;
          intData2acc_RNIBRV9_1               : out   std_logic;
          intData2acc_RNIBRV9_3               : out   std_logic;
          Main_ctl4SD_0_ByteRdEn              : out   std_logic;
          CMOS_DrvX_0_LVDSen_1                : in    std_logic;
          CMOS_DrvX_0_LVDSen_2                : in    std_logic;
          Main_ctl4SD_0_Fifo_wr               : out   std_logic;
          Main_ctl4SD_0_fifo_rd               : out   std_logic;
          \Z\\Fifo_rd_0_Q_[71]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[70]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[69]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[68]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[67]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[66]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[65]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[64]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[63]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[62]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[61]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[60]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[59]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[58]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[57]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[56]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[55]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[54]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[53]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[52]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[51]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[50]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[49]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[48]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[47]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[46]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[45]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[44]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[43]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[42]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[41]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[40]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[39]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[38]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[37]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[36]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[35]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[34]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[33]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[32]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[31]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[30]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[29]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[28]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[27]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[26]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[25]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[24]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[23]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[22]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[21]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[20]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[19]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[18]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[17]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[16]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[15]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[14]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[13]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[12]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[11]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[10]\\\             : in    std_logic;
          \Z\\Fifo_rd_0_Q_[9]\\\              : in    std_logic;
          \Z\\Fifo_rd_0_Q_[8]\\\              : in    std_logic;
          \Z\\Fifo_rd_0_Q_[7]\\\              : in    std_logic;
          \Z\\Fifo_rd_0_Q_[6]\\\              : in    std_logic;
          \Z\\Fifo_rd_0_Q_[5]\\\              : in    std_logic;
          \Z\\Fifo_rd_0_Q_[4]\\\              : in    std_logic;
          \Z\\Fifo_rd_0_Q_[3]\\\              : in    std_logic;
          \Z\\Fifo_rd_0_Q_[2]\\\              : in    std_logic;
          \Z\\Fifo_rd_0_Q_[1]\\\              : in    std_logic;
          \Z\\Fifo_rd_0_Q_[0]\\\              : in    std_logic;
          CMOS_DrvX_0_SDramEn_2               : in    std_logic;
          CMOS_DrvX_0_SDramEn_1               : in    std_logic;
          CMOS_DrvX_0_SDramEn                 : in    std_logic;
          CMOS_DrvX_0_SDramEn_5               : in    std_logic;
          CMOS_DrvX_0_SDramEn_4               : in    std_logic;
          CMOS_DrvX_0_SDramEn_3               : in    std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[71]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[70]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[69]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[68]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[67]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[66]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[65]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[64]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[63]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[62]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[61]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[60]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[59]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[58]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[57]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[56]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[55]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[54]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[53]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[52]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[51]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[50]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[49]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[48]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[47]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[46]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[45]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[44]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[43]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[42]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[41]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[40]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[39]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[38]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[37]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[36]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[35]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[34]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[33]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[32]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[31]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[30]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[29]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[28]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[27]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[26]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[25]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[24]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[23]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[22]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[21]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[20]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[19]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[18]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[17]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[16]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[15]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[14]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[13]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[12]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[11]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[10]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[9]\\\  : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[8]\\\  : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[7]\\\  : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[6]\\\  : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[5]\\\  : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[4]\\\  : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[3]\\\  : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[2]\\\  : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[1]\\\  : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[0]\\\  : out   std_logic;
          Main_ctl4SD_0_fifo_rst_n            : out   std_logic;
          FrameMk_0_LVDS_ok                   : in    std_logic;
          CMOS_DrvX_0_SDramEn_0               : in    std_logic;
          LVDS_enReg                          : in    std_logic;
          un6_sdramenreg                      : out   std_logic;
          CMOS_DrvX_0_AdcEn                   : in    std_logic;
          N_6                                 : out   std_logic;
          N_4                                 : out   std_logic;
          \Z\\My_adder0_0_Sum_[3]\\\          : in    std_logic;
          \Z\\My_adder0_0_Sum_[2]\\\          : in    std_logic;
          \Z\\My_adder0_0_Sum_[1]\\\          : in    std_logic;
          \Z\\My_adder0_0_Sum_[0]\\\          : in    std_logic;
          \Z\\My_adder0_0_Sum_[7]\\\          : in    std_logic;
          \Z\\My_adder0_0_Sum_[6]\\\          : in    std_logic;
          \Z\\My_adder0_0_Sum_[5]\\\          : in    std_logic;
          \Z\\My_adder0_0_Sum_[4]\\\          : in    std_logic;
          \Z\\My_adder0_0_Sum_[11]\\\         : in    std_logic;
          \Z\\My_adder0_0_Sum_[10]\\\         : in    std_logic;
          \Z\\My_adder0_0_Sum_[9]\\\          : in    std_logic;
          \Z\\My_adder0_0_Sum_[8]\\\          : in    std_logic;
          \Z\\My_adder0_0_Sum_[15]\\\         : in    std_logic;
          \Z\\My_adder0_0_Sum_[14]\\\         : in    std_logic;
          \Z\\My_adder0_0_Sum_[13]\\\         : in    std_logic;
          \Z\\My_adder0_0_Sum_[12]\\\         : in    std_logic;
          \Z\\My_adder0_2_Sum_[1]\\\          : in    std_logic;
          \Z\\My_adder0_2_Sum_[0]\\\          : in    std_logic;
          \Z\\My_adder0_1_Sum_[8]\\\          : in    std_logic;
          \Z\\My_adder0_0_Sum_[16]\\\         : in    std_logic;
          \Z\\My_adder0_2_Sum_[3]\\\          : in    std_logic;
          \Z\\My_adder0_2_Sum_[2]\\\          : in    std_logic;
          \Z\\My_adder0_1_Sum_[9]\\\          : in    std_logic;
          \Z\\My_adder0_0_Sum_[17]\\\         : in    std_logic;
          \Z\\My_adder0_2_Sum_[5]\\\          : in    std_logic;
          \Z\\My_adder0_2_Sum_[4]\\\          : in    std_logic;
          \Z\\My_adder0_1_Sum_[10]\\\         : in    std_logic;
          \Z\\My_adder0_1_Sum_[0]\\\          : in    std_logic;
          \Z\\My_adder0_2_Sum_[7]\\\          : in    std_logic;
          \Z\\My_adder0_2_Sum_[6]\\\          : in    std_logic;
          \Z\\My_adder0_1_Sum_[11]\\\         : in    std_logic;
          \Z\\My_adder0_1_Sum_[1]\\\          : in    std_logic;
          \Z\\My_adder0_2_Sum_[9]\\\          : in    std_logic;
          \Z\\My_adder0_2_Sum_[8]\\\          : in    std_logic;
          \Z\\My_adder0_1_Sum_[12]\\\         : in    std_logic;
          \Z\\My_adder0_1_Sum_[2]\\\          : in    std_logic;
          \Z\\My_adder0_2_Sum_[11]\\\         : in    std_logic;
          \Z\\My_adder0_2_Sum_[10]\\\         : in    std_logic;
          \Z\\My_adder0_1_Sum_[13]\\\         : in    std_logic;
          \Z\\My_adder0_1_Sum_[3]\\\          : in    std_logic;
          \Z\\My_adder0_2_Sum_[13]\\\         : in    std_logic;
          \Z\\My_adder0_2_Sum_[12]\\\         : in    std_logic;
          \Z\\My_adder0_1_Sum_[14]\\\         : in    std_logic;
          \Z\\My_adder0_1_Sum_[4]\\\          : in    std_logic;
          \Z\\My_adder0_2_Sum_[15]\\\         : in    std_logic;
          \Z\\My_adder0_2_Sum_[14]\\\         : in    std_logic;
          \Z\\My_adder0_1_Sum_[15]\\\         : in    std_logic;
          \Z\\My_adder0_1_Sum_[5]\\\          : in    std_logic;
          \Z\\My_adder0_2_Sum_[17]\\\         : in    std_logic;
          \Z\\My_adder0_2_Sum_[16]\\\         : in    std_logic;
          \Z\\My_adder0_1_Sum_[16]\\\         : in    std_logic;
          \Z\\My_adder0_1_Sum_[6]\\\          : in    std_logic;
          \Z\\My_adder0_3_Sum_[1]\\\          : in    std_logic;
          \Z\\My_adder0_3_Sum_[0]\\\          : in    std_logic;
          \Z\\My_adder0_1_Sum_[17]\\\         : in    std_logic;
          \Z\\My_adder0_1_Sum_[7]\\\          : in    std_logic;
          \Z\\My_adder0_3_Sum_[5]\\\          : in    std_logic;
          \Z\\My_adder0_3_Sum_[4]\\\          : in    std_logic;
          \Z\\My_adder0_3_Sum_[3]\\\          : in    std_logic;
          \Z\\My_adder0_3_Sum_[2]\\\          : in    std_logic;
          \Z\\My_adder0_3_Sum_[9]\\\          : in    std_logic;
          \Z\\My_adder0_3_Sum_[8]\\\          : in    std_logic;
          \Z\\My_adder0_3_Sum_[7]\\\          : in    std_logic;
          \Z\\My_adder0_3_Sum_[6]\\\          : in    std_logic;
          \Z\\My_adder0_3_Sum_[13]\\\         : in    std_logic;
          \Z\\My_adder0_3_Sum_[12]\\\         : in    std_logic;
          \Z\\My_adder0_3_Sum_[11]\\\         : in    std_logic;
          \Z\\My_adder0_3_Sum_[10]\\\         : in    std_logic;
          \Z\\My_adder0_3_Sum_[17]\\\         : in    std_logic;
          \Z\\My_adder0_3_Sum_[16]\\\         : in    std_logic;
          \Z\\My_adder0_3_Sum_[15]\\\         : in    std_logic;
          \Z\\My_adder0_3_Sum_[14]\\\         : in    std_logic;
          FrameMk_0_LVDS_ok_i                 : in    std_logic;
          Main_ctl4SD_0_fifo_rst_n_0          : out   std_logic;
          Main_ctl4SD_0_fifo_rst_n_1          : out   std_logic;
          Main_ctl4SD_0_fifo_rst_n_2          : out   std_logic;
          Main_ctl4SD_0_fifo_rst_n_3          : out   std_logic;
          Main_ctl4SD_0_fifo_rst_n_4          : out   std_logic;
          Main_ctl4SD_0_fifo_rst_n_5          : out   std_logic;
          PLL_Test1_0_SysRst_O                : in    std_logic;
          PLL_Test1_0_Sys_66M_Clk             : in    std_logic;
          Main_ctl4SD_0_fifo_rst_n_6          : out   std_logic
        );

end Main_ctl4SD;

architecture DEF_ARCH of Main_ctl4SD is 

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E0C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component WaveGenSingleZ11
    port( CMOS_DrvX_0_LVDSen_2    : in    std_logic := 'U';
          CMOS_DrvX_0_LVDSen_1    : in    std_logic := 'U';
          lvdsFifoRowRdOut        : out   std_logic;
          lvdsFifoRowRdOut_i      : out   std_logic;
          PLL_Test1_0_SysRst_O    : in    std_logic := 'U';
          PLL_Test1_0_Sys_66M_Clk : in    std_logic := 'U'
        );
  end component;

  component WaveGenSingleZ14
    port( PrState_2               : in    std_logic := 'U';
          PrState_0               : in    std_logic_vector(4 to 4) := (others => 'U');
          PLL_Test1_0_SysRst_O    : in    std_logic := 'U';
          PLL_Test1_0_Sys_66M_Clk : in    std_logic := 'U';
          latch4acc_0_sqmuxa      : out   std_logic;
          FifoRowRdOut_1          : in    std_logic := 'U';
          FifoRowRdOut_0          : in    std_logic := 'U';
          latch4acc_0_sqmuxa_0    : out   std_logic;
          CMOS_DrvX_0_SDramEn_0   : in    std_logic := 'U';
          latch4acc_0_sqmuxa_1    : out   std_logic
        );
  end component;

  component WaveGenSingleZ8
    port( lvdsFifoRowRdOut_i      : in    std_logic := 'U';
          Main_ctl4SD_0_ByteRdEn  : out   std_logic;
          PLL_Test1_0_SysRst_O    : in    std_logic := 'U';
          PLL_Test1_0_Sys_66M_Clk : in    std_logic := 'U';
          lvdsFifoRowRdOut        : in    std_logic := 'U'
        );
  end component;

  component WaveGenSingleZ12
    port( PrState_4               : out   std_logic;
          PrState_0               : out   std_logic_vector(4 to 4);
          latch_en                : out   std_logic;
          FifoRowRdOut            : in    std_logic := 'U';
          FifoRowRdOut_0          : in    std_logic := 'U';
          PLL_Test1_0_SysRst_O    : in    std_logic := 'U';
          FifoRowRdOut_i          : in    std_logic := 'U';
          PLL_Test1_0_Sys_66M_Clk : in    std_logic := 'U'
        );
  end component;

  component WaveGenSingleZ16
    port( PrState_2               : in    std_logic := 'U';
          PrState_0               : in    std_logic_vector(4 to 4) := (others => 'U');
          PLL_Test1_0_SysRst_O    : in    std_logic := 'U';
          PLL_Test1_0_Sys_66M_Clk : in    std_logic := 'U';
          lvds_fifoRd             : in    std_logic := 'U';
          Main_ctl4SD_0_fifo_rd   : out   std_logic;
          FifoRowRdOut_1          : in    std_logic := 'U';
          FifoRowRdOut_0          : in    std_logic := 'U'
        );
  end component;

  component WaveGenSingleZ17
    port( FifoRowRdOut            : out   std_logic;
          CMOS_DrvX_0_SDramEn_0   : in    std_logic := 'U';
          FifoRowRdOut_i          : out   std_logic;
          FifoRowRdOut_0          : out   std_logic;
          FifoRowRdOut_1          : out   std_logic;
          PLL_Test1_0_SysRst_O    : in    std_logic := 'U';
          PLL_Test1_0_Sys_66M_Clk : in    std_logic := 'U';
          FifoRowRdOut_2          : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component WaveGenSingleZ10
    port( lvds_fifoRd             : out   std_logic;
          PLL_Test1_0_SysRst_O    : in    std_logic := 'U';
          PLL_Test1_0_Sys_66M_Clk : in    std_logic := 'U';
          lvdsFifoRowRdOut        : in    std_logic := 'U'
        );
  end component;

  component WaveGenSingleZ15
    port( Main_ctl4SD_0_Fifo_wr   : out   std_logic;
          PLL_Test1_0_SysRst_O    : in    std_logic := 'U';
          PLL_Test1_0_Sys_66M_Clk : in    std_logic := 'U';
          FifoRowRdOut_1          : in    std_logic := 'U';
          FifoRowRdOut_0          : in    std_logic := 'U'
        );
  end component;

  component WaveGenSingleZ13
    port( PLL_Test1_0_SysRst_O    : in    std_logic := 'U';
          PLL_Test1_0_Sys_66M_Clk : in    std_logic := 'U';
          FifoRowRdOut            : in    std_logic := 'U';
          Data2Fifo_0_sqmuxa      : out   std_logic;
          FifoRowRdOut_1          : in    std_logic := 'U';
          FifoRowRdOut_0          : in    std_logic := 'U';
          Data2Fifo_0_sqmuxa_0    : out   std_logic;
          CMOS_DrvX_0_SDramEn_0   : in    std_logic := 'U';
          Data2Fifo_0_sqmuxa_1    : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \notfirstFrame_0\, \intData2acc[55]_net_1\, 
        FifoRowRdOut_0, \intData2acc[54]_net_1\, 
        \notfirstFrame_1\, \notfirstFrame_1_sqmuxa\, 
        \intData2acc[20]_net_1\, \intData2acc[2]_net_1\, 
        \intData2acc[37]_net_1\, \intData2acc[19]_net_1\, 
        \intData2acc[1]_net_1\, \intData2acc[36]_net_1\, 
        \intData2acc[18]_net_1\, \intData2acc[0]_net_1\, N_8, 
        \latch_data[68]_net_1\, N_15, N_10, 
        \latch_data[69]_net_1\, N_12, \latch_data[70]_net_1\, 
        N_14, \latch_data[71]_net_1\, N_1348, 
        \latch_data[64]_net_1\, N_1349, \latch_data[65]_net_1\, 
        N_1350, \latch_data[66]_net_1\, N_1351, 
        \latch_data[67]_net_1\, N_1367, \latch_data[60]_net_1\, 
        N_1368, \latch_data[61]_net_1\, N_1369, 
        \latch_data[62]_net_1\, N_1370, \latch_data[63]_net_1\, 
        N_1386, \latch_data[56]_net_1\, N_1387, 
        \latch_data[57]_net_1\, N_1388, \latch_data[58]_net_1\, 
        N_1389, \latch_data[59]_net_1\, N_1405, 
        \latch_data[25]_net_1\, N_1546, N_1406, 
        \latch_data[35]_net_1\, N_1407, \latch_data[54]_net_1\, 
        N_1408, \latch_data[55]_net_1\, \ChSel[1]_net_1\, 
        \ChSel[0]_net_1\, N_1422, \latch_data[24]_net_1\, N_1423, 
        \latch_data[34]_net_1\, N_1424, \latch_data[52]_net_1\, 
        N_1585, N_1425, \latch_data[53]_net_1\, N_1442, 
        \latch_data[23]_net_1\, N_1443, \latch_data[33]_net_1\, 
        N_1444, \latch_data[50]_net_1\, N_1445, 
        \latch_data[51]_net_1\, N_1462, \latch_data[22]_net_1\, 
        N_1463, \latch_data[32]_net_1\, N_1464, 
        \latch_data[48]_net_1\, N_1465, \latch_data[49]_net_1\, 
        N_1482, \latch_data[21]_net_1\, N_1483, 
        \latch_data[31]_net_1\, N_1484, \latch_data[46]_net_1\, 
        N_1485, \latch_data[47]_net_1\, N_1502, 
        \latch_data[20]_net_1\, N_1503, \latch_data[30]_net_1\, 
        N_1504, \latch_data[44]_net_1\, N_1505, 
        \latch_data[45]_net_1\, N_1522, \latch_data[19]_net_1\, 
        N_1523, \latch_data[29]_net_1\, N_1524, 
        \latch_data[42]_net_1\, N_1525, \latch_data[43]_net_1\, 
        N_1542, \latch_data[18]_net_1\, N_1543, 
        \latch_data[28]_net_1\, N_1544, \latch_data[40]_net_1\, 
        N_1545, \latch_data[41]_net_1\, N_1562, 
        \latch_data[17]_net_1\, N_1657, N_1563, 
        \latch_data[27]_net_1\, N_1564, \latch_data[38]_net_1\, 
        N_1565, \latch_data[39]_net_1\, N_1581, 
        \latch_data[16]_net_1\, N_1582, \latch_data[26]_net_1\, 
        N_1583, \latch_data[36]_net_1\, N_1584, 
        \latch_data[37]_net_1\, N_1602, \latch_data[12]_net_1\, 
        N_1603, \latch_data[13]_net_1\, N_1604, 
        \latch_data[14]_net_1\, N_1605, \latch_data[15]_net_1\, 
        N_1619, \latch_data[8]_net_1\, N_1620, 
        \latch_data[9]_net_1\, N_1621, \latch_data[10]_net_1\, 
        N_1622, \latch_data[11]_net_1\, N_1636, 
        \latch_data[4]_net_1\, N_1637, \latch_data[5]_net_1\, 
        N_1638, \latch_data[6]_net_1\, N_1639, 
        \latch_data[7]_net_1\, N_1653, \latch_data[0]_net_1\, 
        N_1654, \latch_data[1]_net_1\, N_1655, 
        \latch_data[2]_net_1\, N_1656, \latch_data[3]_net_1\, 
        FifoRowRdOut_1, \intData2acc[68]_net_1\, 
        \intData2acc[69]_net_1\, \intData2acc[70]_net_1\, N_1671, 
        \latch4acc[68]_net_1\, N_1766, N_1672, 
        \latch4acc[69]_net_1\, N_1673, \latch4acc[70]_net_1\, 
        \intData2acc[65]_net_1\, \intData2acc[66]_net_1\, 
        \intData2acc[67]_net_1\, N_1687, \latch4acc[65]_net_1\, 
        N_1688, \latch4acc[66]_net_1\, N_1689, 
        \latch4acc[67]_net_1\, \intData2acc[62]_net_1\, 
        \intData2acc[63]_net_1\, \intData2acc[64]_net_1\, N_1706, 
        \latch4acc[62]_net_1\, N_1707, \latch4acc[63]_net_1\, 
        N_1708, \latch4acc[64]_net_1\, \intData2acc[59]_net_1\, 
        \intData2acc[60]_net_1\, \intData2acc[61]_net_1\, N_1725, 
        \latch4acc[59]_net_1\, N_1726, \latch4acc[60]_net_1\, 
        N_1727, \latch4acc[61]_net_1\, \intData2acc[56]_net_1\, 
        \intData2acc[57]_net_1\, \intData2acc[58]_net_1\, N_1744, 
        \latch4acc[56]_net_1\, N_1745, \latch4acc[57]_net_1\, 
        N_1746, \latch4acc[58]_net_1\, \intData2acc[53]_net_1\, 
        N_1763, \latch4acc[53]_net_1\, N_1876, N_1764, 
        \latch4acc[54]_net_1\, N_1765, \latch4acc[55]_net_1\, 
        \addSel[1]_net_1\, \addSel[0]_net_1\, 
        \intData2acc[50]_net_1\, \intData2acc[51]_net_1\, 
        FifoRowRdOut_2, \intData2acc[52]_net_1\, N_1783, 
        \latch4acc[50]_net_1\, N_1784, \latch4acc[51]_net_1\, 
        N_1785, \latch4acc[52]_net_1\, \intData2acc[47]_net_1\, 
        \intData2acc[48]_net_1\, \intData2acc[49]_net_1\, N_1801, 
        \latch4acc[47]_net_1\, N_1802, \latch4acc[48]_net_1\, 
        N_1803, \latch4acc[49]_net_1\, \intData2acc[44]_net_1\, 
        \intData2acc[45]_net_1\, \intData2acc[46]_net_1\, N_1819, 
        \latch4acc[44]_net_1\, N_1820, \latch4acc[45]_net_1\, 
        N_1821, \latch4acc[46]_net_1\, \intData2acc[41]_net_1\, 
        \intData2acc[42]_net_1\, \intData2acc[43]_net_1\, N_1837, 
        \latch4acc[41]_net_1\, N_1838, \latch4acc[42]_net_1\, 
        N_1839, \latch4acc[43]_net_1\, \intData2acc[38]_net_1\, 
        \intData2acc[39]_net_1\, \intData2acc[40]_net_1\, N_1855, 
        \latch4acc[38]_net_1\, N_1856, \latch4acc[39]_net_1\, 
        N_1857, \latch4acc[40]_net_1\, \intData2acc[35]_net_1\, 
        N_1873, \latch4acc[35]_net_1\, N_1986, N_1874, 
        \latch4acc[36]_net_1\, N_1875, \latch4acc[37]_net_1\, 
        \intData2acc[32]_net_1\, \intData2acc[33]_net_1\, 
        \intData2acc[34]_net_1\, N_1893, \latch4acc[32]_net_1\, 
        N_1894, \latch4acc[33]_net_1\, N_1895, 
        \latch4acc[34]_net_1\, \intData2acc[29]_net_1\, 
        \intData2acc[30]_net_1\, \intData2acc[31]_net_1\, N_1911, 
        \latch4acc[29]_net_1\, N_1912, \latch4acc[30]_net_1\, 
        N_1913, \latch4acc[31]_net_1\, \notfirstFrame\, 
        \intData2acc[26]_net_1\, \intData2acc[27]_net_1\, 
        \intData2acc[28]_net_1\, N_1929, \latch4acc[26]_net_1\, 
        N_1930, \latch4acc[27]_net_1\, N_1931, 
        \latch4acc[28]_net_1\, \intData2acc[23]_net_1\, 
        FifoRowRdOut, \intData2acc[24]_net_1\, 
        \intData2acc[25]_net_1\, N_1947, \latch4acc[23]_net_1\, 
        N_1948, \latch4acc[24]_net_1\, N_1949, 
        \latch4acc[25]_net_1\, \intData2acc[21]_net_1\, 
        \intData2acc[22]_net_1\, N_1965, \latch4acc[20]_net_1\, 
        N_1966, \latch4acc[21]_net_1\, N_1967, 
        \latch4acc[22]_net_1\, \intData2acc[17]_net_1\, N_1983, 
        \latch4acc[17]_net_1\, N_2090, N_1984, 
        \latch4acc[18]_net_1\, N_1985, \latch4acc[19]_net_1\, 
        \intData2acc[14]_net_1\, \intData2acc[15]_net_1\, 
        \intData2acc[16]_net_1\, N_2002, \latch4acc[14]_net_1\, 
        N_2003, \latch4acc[15]_net_1\, N_2004, 
        \latch4acc[16]_net_1\, \intData2acc[11]_net_1\, 
        \intData2acc[12]_net_1\, \intData2acc[13]_net_1\, N_2019, 
        \latch4acc[11]_net_1\, N_2020, \latch4acc[12]_net_1\, 
        N_2021, \latch4acc[13]_net_1\, \intData2acc[8]_net_1\, 
        \intData2acc[9]_net_1\, \intData2acc[10]_net_1\, N_2036, 
        \latch4acc[8]_net_1\, N_2037, \latch4acc[9]_net_1\, 
        N_2038, \latch4acc[10]_net_1\, \intData2acc[5]_net_1\, 
        \intData2acc[6]_net_1\, \intData2acc[7]_net_1\, N_2053, 
        \latch4acc[5]_net_1\, N_2054, \latch4acc[6]_net_1\, 
        N_2055, \latch4acc[7]_net_1\, \intData2acc[3]_net_1\, 
        \intData2acc[4]_net_1\, N_2070, \latch4acc[2]_net_1\, 
        N_2071, \latch4acc[3]_net_1\, N_2072, 
        \latch4acc[4]_net_1\, \ChSel_3[0]\, latch_en, 
        \ChSel_3[1]\, \addSel_2[0]\, \addSel_2[1]\, 
        \intData2acc[71]_net_1\, N_2087, \latch4acc[0]_net_1\, 
        N_2088, \latch4acc[1]_net_1\, N_2089, 
        \latch4acc[71]_net_1\, un6_sdramenreg_net_1, 
        Data2Fifo_0_sqmuxa_0, Data2Fifo_0_sqmuxa_1, 
        Data2Fifo_0_sqmuxa, latch4acc_0_sqmuxa_0, 
        latch4acc_0_sqmuxa_1, latch4acc_0_sqmuxa, FifoRowRdOut_i, 
        \PrState[4]\, \PrState_0[4]\, lvds_fifoRd, 
        lvdsFifoRowRdOut, lvdsFifoRowRdOut_i, \GND\, \VCC\, GND_0, 
        VCC_0 : std_logic;

    for all : WaveGenSingleZ11
	Use entity work.WaveGenSingleZ11(DEF_ARCH);
    for all : WaveGenSingleZ14
	Use entity work.WaveGenSingleZ14(DEF_ARCH);
    for all : WaveGenSingleZ8
	Use entity work.WaveGenSingleZ8(DEF_ARCH);
    for all : WaveGenSingleZ12
	Use entity work.WaveGenSingleZ12(DEF_ARCH);
    for all : WaveGenSingleZ16
	Use entity work.WaveGenSingleZ16(DEF_ARCH);
    for all : WaveGenSingleZ17
	Use entity work.WaveGenSingleZ17(DEF_ARCH);
    for all : WaveGenSingleZ10
	Use entity work.WaveGenSingleZ10(DEF_ARCH);
    for all : WaveGenSingleZ15
	Use entity work.WaveGenSingleZ15(DEF_ARCH);
    for all : WaveGenSingleZ13
	Use entity work.WaveGenSingleZ13(DEF_ARCH);
begin 

    un6_sdramenreg <= un6_sdramenreg_net_1;

    \intData2acc_RNI7JV9[34]\ : NOR3C
      port map(A => FifoRowRdOut_2, B => \notfirstFrame_1\, C => 
        \intData2acc[34]_net_1\, Y => intData2acc_RNI7JV9_0);
    
    \intData2acc[35]\ : DFN1E1C0
      port map(D => N_1873, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_1, Q
         => \intData2acc[35]_net_1\);
    
    \intData2acc[20]\ : DFN1E1C0
      port map(D => N_1965, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_1, Q
         => \intData2acc[20]_net_1\);
    
    \latch4acc[45]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[45]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa_1, Q => \latch4acc[45]_net_1\);
    
    \intData2acc_RNIBJV9[38]\ : NOR3C
      port map(A => FifoRowRdOut_2, B => \notfirstFrame_1\, C => 
        \intData2acc[38]_net_1\, Y => intData2acc_RNIBJV9(38));
    
    \intData2acc[21]\ : DFN1E1C0
      port map(D => N_1966, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_1, Q
         => \intData2acc[21]_net_1\);
    
    \latch_data_RNO[9]\ : MX2
      port map(A => \latch_data[9]_net_1\, B => 
        \Z\\My_adder0_0_Sum_[9]\\\, S => N_1657, Y => N_1620);
    
    \latch4acc[44]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[44]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa_1, Q => \latch4acc[44]_net_1\);
    
    notfirstFrame_1 : DFN1E0C0
      port map(D => FrameMk_0_LVDS_ok_i, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => \notfirstFrame_1_sqmuxa\, Q => \notfirstFrame_1\);
    
    \intData2acc_RNICVV9[62]\ : NOR3C
      port map(A => FifoRowRdOut_1, B => \notfirstFrame_0\, C => 
        \intData2acc[62]_net_1\, Y => intData2acc_RNICVV9(62));
    
    \Data2Fifo[61]\ : DFN1E1C0
      port map(D => \latch_data[61]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[61]\\\);
    
    \latch4acc[43]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[43]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa_1, Q => \latch4acc[43]_net_1\);
    
    \latch4acc[41]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[41]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa_1, Q => \latch4acc[41]_net_1\);
    
    \intData2acc_RNIDN36[24]\ : NOR3C
      port map(A => FifoRowRdOut, B => \notfirstFrame\, C => 
        \intData2acc[24]_net_1\, Y => intData2acc_RNIDN36(24));
    
    \latch4acc[56]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[56]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa, Q => \latch4acc[56]_net_1\);
    
    \latch4acc[25]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[25]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa_0, Q => \latch4acc[25]_net_1\);
    
    \intData2acc_RNICNV9[46]\ : NOR3C
      port map(A => FifoRowRdOut_2, B => \notfirstFrame_1\, C => 
        \intData2acc[46]_net_1\, Y => intData2acc_RNICNV9(46));
    
    \latch_data_RNO[3]\ : MX2
      port map(A => \latch_data[3]_net_1\, B => 
        \Z\\My_adder0_0_Sum_[3]\\\, S => N_1657, Y => N_1656);
    
    \latch_data[9]\ : DFN1E1C0
      port map(D => N_1620, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn, Q => 
        \latch_data[9]_net_1\);
    
    \latch4acc[24]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[24]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa_0, Q => \latch4acc[24]_net_1\);
    
    \intData2acc_RNI0KS7[26]\ : NOR3C
      port map(A => FifoRowRdOut_2, B => \notfirstFrame\, C => 
        \intData2acc[26]_net_1\, Y => intData2acc_RNI0KS7(26));
    
    \intData2acc[6]\ : DFN1E1C0
      port map(D => N_2054, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_3, Q
         => \intData2acc[6]_net_1\);
    
    \latch4acc[23]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[23]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa_0, Q => \latch4acc[23]_net_1\);
    
    \latch4acc[21]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[21]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa_0, Q => \latch4acc[21]_net_1\);
    
    \latch4acc[68]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[68]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa, Q => \latch4acc[68]_net_1\);
    
    \intData2acc_RNI5JV9[32]\ : NOR3C
      port map(A => FifoRowRdOut_2, B => \notfirstFrame_1\, C => 
        \intData2acc[32]_net_1\, Y => intData2acc_RNI5JV9(32));
    
    \latch4acc[50]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[50]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa_1, Q => \latch4acc[50]_net_1\);
    
    \intData2acc[58]\ : DFN1E1C0
      port map(D => N_1746, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_3, Q
         => \intData2acc[58]_net_1\);
    
    \Data2Fifo[12]\ : DFN1E1C0
      port map(D => \latch_data[12]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa_0, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[12]\\\);
    
    \Data2Fifo[43]\ : DFN1E1C0
      port map(D => \latch_data[43]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa_1, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[43]\\\);
    
    \Data2Fifo[20]\ : DFN1E1C0
      port map(D => \latch_data[20]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa_0, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[20]\\\);
    
    \latch_data[71]\ : DFN1E1C0
      port map(D => N_14, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn, Q => 
        \latch_data[71]_net_1\);
    
    \intData2acc_RNITJS7[23]\ : NOR3C
      port map(A => FifoRowRdOut_2, B => \notfirstFrame\, C => 
        \intData2acc[23]_net_1\, Y => intData2acc_RNITJS7(23));
    
    \intData2acc_RNIBJ36[15]\ : NOR3C
      port map(A => FifoRowRdOut, B => \notfirstFrame\, C => 
        \intData2acc[15]_net_1\, Y => intData2acc_RNIBJ36(15));
    
    \Data2Fifo[4]\ : DFN1E1C0
      port map(D => \latch_data[4]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa_1, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[4]\\\);
    
    \latch_data[3]\ : DFN1E1C0
      port map(D => N_1656, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_5, Q
         => \latch_data[3]_net_1\);
    
    \latch_data_RNO[71]\ : MX2
      port map(A => \Z\\My_adder0_3_Sum_[17]\\\, B => 
        \latch_data[71]_net_1\, S => N_15, Y => N_14);
    
    \intData2acc[3]\ : DFN1E1C0
      port map(D => N_2071, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_2, Q
         => \intData2acc[3]_net_1\);
    
    \intData2acc_RNO[9]\ : MX2
      port map(A => \latch4acc[9]_net_1\, B => 
        \intData2acc[9]_net_1\, S => N_2090, Y => N_2037);
    
    \latch_data[57]\ : DFN1E1C0
      port map(D => N_1387, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn, Q => 
        \latch_data[57]_net_1\);
    
    \latch4acc[17]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[17]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa_0, Q => \latch4acc[17]_net_1\);
    
    \intData2acc_RNO[1]\ : MX2
      port map(A => \latch4acc[1]_net_1\, B => 
        \intData2acc[1]_net_1\, S => N_2090, Y => N_2088);
    
    \latch_data[36]\ : DFN1E1C0
      port map(D => N_1583, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_5, Q
         => \latch_data[36]_net_1\);
    
    \intData2acc[19]\ : DFN1E1C0
      port map(D => N_1985, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_1, Q
         => \intData2acc[19]_net_1\);
    
    \latch_data_RNO[67]\ : MX2
      port map(A => \Z\\My_adder0_3_Sum_[13]\\\, B => 
        \latch_data[67]_net_1\, S => N_15, Y => N_1351);
    
    \latch_data_RNO[20]\ : MX2
      port map(A => \latch_data[20]_net_1\, B => 
        \Z\\My_adder0_1_Sum_[2]\\\, S => N_1546, Y => N_1502);
    
    \intData2acc_RNO[50]\ : MX2
      port map(A => \latch4acc[50]_net_1\, B => 
        \intData2acc[50]_net_1\, S => N_1876, Y => N_1783);
    
    \Data2Fifo[6]\ : DFN1E1C0
      port map(D => \latch_data[6]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[6]\\\);
    
    \intData2acc_RNIITV6[7]\ : NOR3C
      port map(A => FifoRowRdOut, B => \notfirstFrame\, C => 
        \intData2acc[7]_net_1\, Y => intData2acc_RNIITV6(7));
    
    \latch_data_RNO[28]\ : MX2
      port map(A => \latch_data[28]_net_1\, B => 
        \Z\\My_adder0_1_Sum_[10]\\\, S => N_1546, Y => N_1543);
    
    \intData2acc[32]\ : DFN1E1C0
      port map(D => N_1893, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_1, Q
         => \intData2acc[32]_net_1\);
    
    \intData2acc[10]\ : DFN1E1C0
      port map(D => N_2038, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_0, Q
         => \intData2acc[10]_net_1\);
    
    \latch_data[34]\ : DFN1E1C0
      port map(D => N_1423, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_5, Q
         => \latch_data[34]_net_1\);
    
    \intData2acc[11]\ : DFN1E1C0
      port map(D => N_2019, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_0, Q
         => \intData2acc[11]_net_1\);
    
    \Data2Fifo[51]\ : DFN1E1C0
      port map(D => \latch_data[51]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa_1, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[51]\\\);
    
    notfirstFrame_0 : DFN1E0C0
      port map(D => FrameMk_0_LVDS_ok_i, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => \notfirstFrame_1_sqmuxa\, Q => \notfirstFrame_0\);
    
    \latch_data[62]\ : DFN1E1C0
      port map(D => N_1369, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn, Q => 
        \latch_data[62]_net_1\);
    
    notfirstFrame : DFN1E0C0
      port map(D => FrameMk_0_LVDS_ok_i, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => \notfirstFrame_1_sqmuxa\, Q => \notfirstFrame\);
    
    \latch_data_RNO[22]\ : MX2
      port map(A => \latch_data[22]_net_1\, B => 
        \Z\\My_adder0_1_Sum_[4]\\\, S => N_1546, Y => N_1462);
    
    \latch4acc[58]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[58]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa, Q => \latch4acc[58]_net_1\);
    
    \intData2acc_RNIDNV9[47]\ : NOR3C
      port map(A => FifoRowRdOut_2, B => \notfirstFrame_1\, C => 
        \intData2acc[47]_net_1\, Y => intData2acc_RNIDNV9(47));
    
    \intData2acc[23]\ : DFN1E1C0
      port map(D => N_1947, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_1, Q
         => \intData2acc[23]_net_1\);
    
    \Data2Fifo[28]\ : DFN1E1C0
      port map(D => \latch_data[28]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa_0, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[28]\\\);
    
    fifo_rst_n_2 : DFN1C0
      port map(D => pr_state_ns(8), CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => Main_ctl4SD_0_fifo_rst_n_2);
    
    \Data2Fifo[46]\ : DFN1E1C0
      port map(D => \latch_data[46]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa_1, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[46]\\\);
    
    \intData2acc_RNO[35]\ : MX2
      port map(A => \latch4acc[35]_net_1\, B => 
        \intData2acc[35]_net_1\, S => N_1986, Y => N_1873);
    
    \intData2acc_RNI4JV9[31]\ : NOR3C
      port map(A => FifoRowRdOut_2, B => \notfirstFrame_1\, C => 
        \intData2acc[31]_net_1\, Y => intData2acc_RNI4JV9(31));
    
    \latch_data_RNO[47]\ : MX2
      port map(A => \Z\\My_adder0_2_Sum_[11]\\\, B => 
        \latch_data[47]_net_1\, S => N_1585, Y => N_1485);
    
    \latch_data_RNO[33]\ : MX2
      port map(A => \latch_data[33]_net_1\, B => 
        \Z\\My_adder0_1_Sum_[15]\\\, S => N_1546, Y => N_1443);
    
    \intData2acc_RNID30A[70]\ : NOR3C
      port map(A => FifoRowRdOut_1, B => \notfirstFrame_0\, C => 
        \intData2acc[70]_net_1\, Y => intData2acc_RNID30A(70));
    
    \addSel_RNO[0]\ : NOR2
      port map(A => \addSel[0]_net_1\, B => CMOS_DrvX_0_AdcEn, Y
         => \addSel_2[0]\);
    
    \latch4acc[32]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[32]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa_1, Q => \latch4acc[32]_net_1\);
    
    \intData2acc[5]\ : DFN1E1C0
      port map(D => N_2053, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_3, Q
         => \intData2acc[5]_net_1\);
    
    \latch4acc[71]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[71]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa, Q => \latch4acc[71]_net_1\);
    
    \intData2acc_RNO[45]\ : MX2
      port map(A => \latch4acc[45]_net_1\, B => 
        \intData2acc[45]_net_1\, S => N_1876, Y => N_1820);
    
    \Data2Fifo[31]\ : DFN1E1C0
      port map(D => \latch_data[31]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa_1, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[31]\\\);
    
    \intData2acc[47]\ : DFN1E1C0
      port map(D => N_1801, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_2, Q
         => \intData2acc[47]_net_1\);
    
    \latch4acc[5]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[5]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa, Q => \latch4acc[5]_net_1\);
    
    \intData2acc_RNO[56]\ : MX2
      port map(A => \latch4acc[56]_net_1\, B => 
        \intData2acc[56]_net_1\, S => N_1766, Y => N_1744);
    
    \intData2acc_RNIBRV9[53]\ : NOR3C
      port map(A => FifoRowRdOut_1, B => \notfirstFrame_1\, C => 
        \intData2acc[53]_net_1\, Y => intData2acc_RNIBRV9_1);
    
    \intData2acc[28]\ : DFN1E1C0
      port map(D => N_1931, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_1, Q
         => \intData2acc[28]_net_1\);
    
    \ChSel_RNITABA_2[1]\ : NOR2
      port map(A => \ChSel[1]_net_1\, B => \ChSel[0]_net_1\, Y
         => N_1657);
    
    \latch_data[43]\ : DFN1E1C0
      port map(D => N_1525, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_5, Q
         => \latch_data[43]_net_1\);
    
    \intData2acc_RNO[22]\ : MX2
      port map(A => \latch4acc[22]_net_1\, B => 
        \intData2acc[22]_net_1\, S => N_1986, Y => N_1967);
    
    \latch_data_RNO[8]\ : MX2
      port map(A => \latch_data[8]_net_1\, B => 
        \Z\\My_adder0_0_Sum_[8]\\\, S => N_1657, Y => N_1619);
    
    \Data2Fifo[24]\ : DFN1E1C0
      port map(D => \latch_data[24]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa_0, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[24]\\\);
    
    \intData2acc[1]\ : DFN1E1C0
      port map(D => N_2088, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_1, Q
         => \intData2acc[1]_net_1\);
    
    \latch_data_RNO[1]\ : MX2
      port map(A => \latch_data[1]_net_1\, B => 
        \Z\\My_adder0_0_Sum_[1]\\\, S => N_1657, Y => N_1654);
    
    \intData2acc[39]\ : DFN1E1C0
      port map(D => N_1856, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_2, Q
         => \intData2acc[39]_net_1\);
    
    \Data2Fifo[5]\ : DFN1E1C0
      port map(D => \latch_data[5]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[5]\\\);
    
    \intData2acc_RNIHVV9[67]\ : NOR3C
      port map(A => FifoRowRdOut_1, B => \notfirstFrame_0\, C => 
        \intData2acc[67]_net_1\, Y => intData2acc_RNIHVV9(67));
    
    \intData2acc[67]\ : DFN1E1C0
      port map(D => N_1689, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_3, Q
         => \intData2acc[67]_net_1\);
    
    \intData2acc[56]\ : DFN1E1C0
      port map(D => N_1744, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_2, Q
         => \intData2acc[56]_net_1\);
    
    \addSel_RNILVIF[1]\ : OR2B
      port map(A => \addSel[1]_net_1\, B => \addSel[0]_net_1\, Y
         => N_1766);
    
    \latch_data[45]\ : DFN1E1C0
      port map(D => N_1505, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_5, Q
         => \latch_data[45]_net_1\);
    
    \latch_data[28]\ : DFN1E1C0
      port map(D => N_1543, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_4, Q
         => \latch_data[28]_net_1\);
    
    \intData2acc_RNIBNV9[45]\ : NOR3C
      port map(A => FifoRowRdOut_2, B => \notfirstFrame_1\, C => 
        \intData2acc[45]_net_1\, Y => intData2acc_RNIBNV9(45));
    
    \latch_data_RNO[14]\ : MX2
      port map(A => \latch_data[14]_net_1\, B => 
        \Z\\My_adder0_0_Sum_[14]\\\, S => N_1657, Y => N_1604);
    
    \intData2acc_RNI3BV9[19]\ : NOR3C
      port map(A => \notfirstFrame_0\, B => 
        \intData2acc[19]_net_1\, C => FifoRowRdOut_0, Y => 
        intData2acc_RNI3BV9(19));
    
    \intData2acc[30]\ : DFN1E1C0
      port map(D => N_1912, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_1, Q
         => \intData2acc[30]_net_1\);
    
    \ChSel_RNITABA_1[1]\ : NOR2A
      port map(A => \ChSel[0]_net_1\, B => \ChSel[1]_net_1\, Y
         => N_1546);
    
    \latch_data[21]\ : DFN1E1C0
      port map(D => N_1482, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_4, Q
         => \latch_data[21]_net_1\);
    
    \intData2acc[13]\ : DFN1E1C0
      port map(D => N_2021, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_0, Q
         => \intData2acc[13]_net_1\);
    
    \intData2acc[31]\ : DFN1E1C0
      port map(D => N_1913, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_1, Q
         => \intData2acc[31]_net_1\);
    
    \latch_data[29]\ : DFN1E1C0
      port map(D => N_1523, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_4, Q
         => \latch_data[29]_net_1\);
    
    fifo_rst_n_4 : DFN1C0
      port map(D => pr_state_ns(8), CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => Main_ctl4SD_0_fifo_rst_n_4);
    
    \intData2acc_RNIEN36[25]\ : NOR3C
      port map(A => FifoRowRdOut, B => \notfirstFrame\, C => 
        \intData2acc[25]_net_1\, Y => intData2acc_RNIEN36(25));
    
    \intData2acc_RNIFNV9[49]\ : NOR3C
      port map(A => FifoRowRdOut_2, B => \notfirstFrame_1\, C => 
        \intData2acc[49]_net_1\, Y => intData2acc_RNIFNV9(49));
    
    \latch_data_RNO[30]\ : MX2
      port map(A => \latch_data[30]_net_1\, B => 
        \Z\\My_adder0_1_Sum_[12]\\\, S => N_1546, Y => N_1503);
    
    \latch_data[56]\ : DFN1E1C0
      port map(D => N_1386, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn, Q => 
        \latch_data[56]_net_1\);
    
    fifo_rst_n_0 : DFN1C0
      port map(D => pr_state_ns(8), CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => Main_ctl4SD_0_fifo_rst_n_0);
    
    \latch_data_RNO[38]\ : MX2
      port map(A => \Z\\My_adder0_2_Sum_[2]\\\, B => 
        \latch_data[38]_net_1\, S => N_1585, Y => N_1564);
    
    \latch_data_RNO[15]\ : MX2
      port map(A => \latch_data[15]_net_1\, B => 
        \Z\\My_adder0_0_Sum_[15]\\\, S => N_1657, Y => N_1605);
    
    \intData2acc_RNO[62]\ : MX2
      port map(A => \latch4acc[62]_net_1\, B => 
        \intData2acc[62]_net_1\, S => N_1766, Y => N_1706);
    
    \intData2acc_RNO[12]\ : MX2
      port map(A => \latch4acc[12]_net_1\, B => 
        \intData2acc[12]_net_1\, S => N_2090, Y => N_2020);
    
    \intData2acc_RNO[51]\ : MX2
      port map(A => \latch4acc[51]_net_1\, B => 
        \intData2acc[51]_net_1\, S => N_1876, Y => N_1784);
    
    \latch_data[54]\ : DFN1E1C0
      port map(D => N_1407, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_5, Q
         => \latch_data[54]_net_1\);
    
    \latch_data_RNO[32]\ : MX2
      port map(A => \latch_data[32]_net_1\, B => 
        \Z\\My_adder0_1_Sum_[14]\\\, S => N_1546, Y => N_1463);
    
    \intData2acc_RNIGVV9[66]\ : NOR3C
      port map(A => FifoRowRdOut_1, B => \notfirstFrame_0\, C => 
        \intData2acc[66]_net_1\, Y => intData2acc_RNIGVV9(66));
    
    \latch4acc[49]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[49]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa_1, Q => \latch4acc[49]_net_1\);
    
    \intData2acc[18]\ : DFN1E1C0
      port map(D => N_1984, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_1, Q
         => \intData2acc[18]_net_1\);
    
    \Data2Fifo[27]\ : DFN1E1C0
      port map(D => \latch_data[27]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa_0, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[27]\\\);
    
    \latch_data_RNO[26]\ : MX2
      port map(A => \latch_data[26]_net_1\, B => 
        \Z\\My_adder0_1_Sum_[8]\\\, S => N_1546, Y => N_1582);
    
    \latch_data[18]\ : DFN1E1C0
      port map(D => N_1542, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_4, Q
         => \latch_data[18]_net_1\);
    
    \intData2acc_RNO[2]\ : MX2
      port map(A => \latch4acc[2]_net_1\, B => 
        \intData2acc[2]_net_1\, S => N_2090, Y => N_2070);
    
    \latch_data_RNO[0]\ : MX2
      port map(A => \latch_data[0]_net_1\, B => 
        \Z\\My_adder0_0_Sum_[0]\\\, S => N_1657, Y => N_1653);
    
    \latch_data[11]\ : DFN1E1C0
      port map(D => N_1622, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_3, Q
         => \latch_data[11]_net_1\);
    
    \latch4acc[36]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[36]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa_1, Q => \latch4acc[36]_net_1\);
    
    \latch4acc[29]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[29]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa_0, Q => \latch4acc[29]_net_1\);
    
    fifo_rst_n : DFN1C0
      port map(D => pr_state_ns(8), CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => Main_ctl4SD_0_fifo_rst_n);
    
    \Data2Fifo[19]\ : DFN1E1C0
      port map(D => \latch_data[19]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa_0, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[19]\\\);
    
    \latch_data[19]\ : DFN1E1C0
      port map(D => N_1522, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_4, Q
         => \latch_data[19]_net_1\);
    
    \ChSel[0]\ : DFN1C0
      port map(D => \ChSel_3[0]\, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \ChSel[0]_net_1\);
    
    \latch_data_RNO[63]\ : MX2
      port map(A => \Z\\My_adder0_3_Sum_[9]\\\, B => 
        \latch_data[63]_net_1\, S => N_15, Y => N_1370);
    
    \latch_data_RNO[6]\ : MX2
      port map(A => \latch_data[6]_net_1\, B => 
        \Z\\My_adder0_0_Sum_[6]\\\, S => N_1657, Y => N_1638);
    
    \latch_data[30]\ : DFN1E1C0
      port map(D => N_1503, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_4, Q
         => \latch_data[30]_net_1\);
    
    \latch4acc[30]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[30]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa_0, Q => \latch4acc[30]_net_1\);
    
    \intData2acc_RNI9J36[13]\ : NOR3C
      port map(A => FifoRowRdOut, B => \notfirstFrame\, C => 
        \intData2acc[13]_net_1\, Y => intData2acc_RNI9J36(13));
    
    \intData2acc_RNI9NV9[43]\ : NOR3C
      port map(A => FifoRowRdOut_2, B => \notfirstFrame_1\, C => 
        \intData2acc[43]_net_1\, Y => intData2acc_RNI9NV9(43));
    
    \latch_data_RNO[19]\ : MX2
      port map(A => \latch_data[19]_net_1\, B => 
        \Z\\My_adder0_1_Sum_[1]\\\, S => N_1546, Y => N_1522);
    
    \latch_data[67]\ : DFN1E1C0
      port map(D => N_1351, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn, Q => 
        \latch_data[67]_net_1\);
    
    \latch_data_RNO[5]\ : MX2
      port map(A => \latch_data[5]_net_1\, B => 
        \Z\\My_adder0_0_Sum_[5]\\\, S => N_1657, Y => N_1637);
    
    \latch4acc[12]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[12]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa_0, Q => \latch4acc[12]_net_1\);
    
    \intData2acc_RNIVOQA[0]\ : NOR3C
      port map(A => \notfirstFrame_0\, B => 
        \intData2acc[0]_net_1\, C => FifoRowRdOut_0, Y => 
        intData2acc_RNIVOQA(0));
    
    \intData2acc[33]\ : DFN1E1C0
      port map(D => N_1894, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_1, Q
         => \intData2acc[33]_net_1\);
    
    \intData2acc[26]\ : DFN1E1C0
      port map(D => N_1929, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_1, Q
         => \intData2acc[26]_net_1\);
    
    \latch_data_RNO[54]\ : MX2
      port map(A => \Z\\My_adder0_3_Sum_[0]\\\, B => 
        \latch_data[54]_net_1\, S => N_15, Y => N_1407);
    
    \intData2acc_RNO[59]\ : MX2
      port map(A => \latch4acc[59]_net_1\, B => 
        \intData2acc[59]_net_1\, S => N_1766, Y => N_1725);
    
    \Data2Fifo[41]\ : DFN1E1C0
      port map(D => \latch_data[41]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa_1, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[41]\\\);
    
    \intData2acc_RNI7J36[11]\ : NOR3C
      port map(A => FifoRowRdOut, B => \notfirstFrame\, C => 
        \intData2acc[11]_net_1\, Y => intData2acc_RNI7J36(11));
    
    \Data2Fifo[60]\ : DFN1E1C0
      port map(D => \latch_data[60]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[60]\\\);
    
    \latch_data_RNO[43]\ : MX2
      port map(A => \Z\\My_adder0_2_Sum_[7]\\\, B => 
        \latch_data[43]_net_1\, S => N_1585, Y => N_1525);
    
    \intData2acc_RNIEVV9[64]\ : NOR3C
      port map(A => FifoRowRdOut_1, B => \notfirstFrame_0\, C => 
        \intData2acc[64]_net_1\, Y => intData2acc_RNIEVV9(64));
    
    \intData2acc_RNO[54]\ : MX2
      port map(A => \latch4acc[54]_net_1\, B => 
        \intData2acc[54]_net_1\, S => N_1766, Y => N_1764);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \latch_data_RNO[55]\ : MX2
      port map(A => \Z\\My_adder0_3_Sum_[1]\\\, B => 
        \latch_data[55]_net_1\, S => N_15, Y => N_1408);
    
    \latch4acc[38]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[38]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa_1, Q => \latch4acc[38]_net_1\);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    \intData2acc_RNO[53]\ : MX2
      port map(A => \latch4acc[53]_net_1\, B => 
        \intData2acc[53]_net_1\, S => N_1876, Y => N_1763);
    
    \intData2acc_RNIBRV9[52]\ : NOR3C
      port map(A => FifoRowRdOut_2, B => \notfirstFrame_1\, C => 
        \intData2acc[52]_net_1\, Y => intData2acc_RNIBRV9_0);
    
    \intData2acc[38]\ : DFN1E1C0
      port map(D => N_1855, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_2, Q
         => \intData2acc[38]_net_1\);
    
    \intData2acc_RNO[57]\ : MX2
      port map(A => \latch4acc[57]_net_1\, B => 
        \intData2acc[57]_net_1\, S => N_1766, Y => N_1745);
    
    \intData2acc_RNIAN36[21]\ : NOR3C
      port map(A => FifoRowRdOut, B => \notfirstFrame\, C => 
        \intData2acc[21]_net_1\, Y => intData2acc_RNIAN36(21));
    
    \Data2Fifo[13]\ : DFN1E1C0
      port map(D => \latch_data[13]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa_0, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[13]\\\);
    
    \addSel[0]\ : DFN1C0
      port map(D => \addSel_2[0]\, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \addSel[0]_net_1\);
    
    \latch_data_RNO[60]\ : MX2
      port map(A => \Z\\My_adder0_3_Sum_[6]\\\, B => 
        \latch_data[60]_net_1\, S => N_15, Y => N_1367);
    
    \intData2acc_RNI7NV9[41]\ : NOR3C
      port map(A => FifoRowRdOut_2, B => \notfirstFrame_1\, C => 
        \intData2acc[41]_net_1\, Y => intData2acc_RNI7NV9(41));
    
    \latch_data_RNO[68]\ : MX2
      port map(A => \Z\\My_adder0_3_Sum_[14]\\\, B => 
        \latch_data[68]_net_1\, S => N_15, Y => N_8);
    
    \intData2acc[8]\ : DFN1E1C0
      port map(D => N_2036, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_3, Q
         => \intData2acc[8]_net_1\);
    
    \Data2Fifo[68]\ : DFN1E1C0
      port map(D => \latch_data[68]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[68]\\\);
    
    \latch_data_RNO[7]\ : MX2
      port map(A => \latch_data[7]_net_1\, B => 
        \Z\\My_adder0_0_Sum_[7]\\\, S => N_1657, Y => N_1639);
    
    \Data2Fifo[25]\ : DFN1E1C0
      port map(D => \latch_data[25]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa_0, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[25]\\\);
    
    \un6_sdramenreg\ : NOR2A
      port map(A => LVDS_enReg, B => CMOS_DrvX_0_SDramEn_0, Y => 
        un6_sdramenreg_net_1);
    
    \latch_data[22]\ : DFN1E1C0
      port map(D => N_1462, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_4, Q
         => \latch_data[22]_net_1\);
    
    \intData2acc_RNIANV9[44]\ : NOR3C
      port map(A => FifoRowRdOut_2, B => \notfirstFrame_1\, C => 
        \intData2acc[44]_net_1\, Y => intData2acc_RNIANV9(44));
    
    \latch_data_RNO[62]\ : MX2
      port map(A => \Z\\My_adder0_3_Sum_[8]\\\, B => 
        \latch_data[62]_net_1\, S => N_15, Y => N_1369);
    
    \latch_data_RNO[36]\ : MX2
      port map(A => \Z\\My_adder0_2_Sum_[0]\\\, B => 
        \latch_data[36]_net_1\, S => N_1585, Y => N_1583);
    
    \intData2acc_RNO[30]\ : MX2
      port map(A => \latch4acc[30]_net_1\, B => 
        \intData2acc[30]_net_1\, S => N_1986, Y => N_1912);
    
    \intData2acc[16]\ : DFN1E1C0
      port map(D => N_2004, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_1, Q
         => \intData2acc[16]_net_1\);
    
    \Data2Fifo[50]\ : DFN1E1C0
      port map(D => \latch_data[50]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa_1, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[50]\\\);
    
    \latch_data_RNO[11]\ : MX2
      port map(A => \latch_data[11]_net_1\, B => 
        \Z\\My_adder0_0_Sum_[11]\\\, S => N_1657, Y => N_1622);
    
    \latch4acc[7]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[7]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa, Q => \latch4acc[7]_net_1\);
    
    \intData2acc_RNO[4]\ : MX2
      port map(A => \latch4acc[4]_net_1\, B => 
        \intData2acc[4]_net_1\, S => N_2090, Y => N_2072);
    
    \latch_data_RNO[59]\ : MX2
      port map(A => \Z\\My_adder0_3_Sum_[5]\\\, B => 
        \latch_data[59]_net_1\, S => N_15, Y => N_1389);
    
    \intData2acc_RNIPB46[71]\ : NOR3C
      port map(A => FifoRowRdOut, B => \notfirstFrame\, C => 
        \intData2acc[71]_net_1\, Y => intData2acc_RNIPB46(71));
    
    \latch4acc[47]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[47]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa_1, Q => \latch4acc[47]_net_1\);
    
    \intData2acc_RNI9RV9[51]\ : NOR3C
      port map(A => FifoRowRdOut_1, B => \notfirstFrame_1\, C => 
        \intData2acc[51]_net_1\, Y => intData2acc_RNI9RV9(51));
    
    \latch_data_RNO[40]\ : MX2
      port map(A => \Z\\My_adder0_2_Sum_[4]\\\, B => 
        \latch_data[40]_net_1\, S => N_1585, Y => N_1544);
    
    \intData2acc_RNO[40]\ : MX2
      port map(A => \latch4acc[40]_net_1\, B => 
        \intData2acc[40]_net_1\, S => N_1876, Y => N_1857);
    
    \intData2acc_RNI6J36[10]\ : NOR3C
      port map(A => FifoRowRdOut, B => \notfirstFrame\, C => 
        \intData2acc[10]_net_1\, Y => intData2acc_RNI6J36(10));
    
    \latch_data_RNO[48]\ : MX2
      port map(A => \Z\\My_adder0_2_Sum_[12]\\\, B => 
        \latch_data[48]_net_1\, S => N_1585, Y => N_1464);
    
    \latch_data[8]\ : DFN1E1C0
      port map(D => N_1619, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn, Q => 
        \latch_data[8]_net_1\);
    
    \latch_data[50]\ : DFN1E1C0
      port map(D => N_1444, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_5, Q
         => \latch_data[50]_net_1\);
    
    \latch4acc[27]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[27]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa_0, Q => \latch4acc[27]_net_1\);
    
    \latch4acc[16]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[16]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa_0, Q => \latch4acc[16]_net_1\);
    
    \Data2Fifo[16]\ : DFN1E1C0
      port map(D => \latch_data[16]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa_0, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[16]\\\);
    
    \latch_data_RNO[42]\ : MX2
      port map(A => \Z\\My_adder0_2_Sum_[6]\\\, B => 
        \latch_data[42]_net_1\, S => N_1585, Y => N_1524);
    
    \intData2acc_RNIBRV9[55]\ : NOR3C
      port map(A => \notfirstFrame_0\, B => 
        \intData2acc[55]_net_1\, C => FifoRowRdOut_0, Y => 
        intData2acc_RNIBRV9_3);
    
    \Data2Fifo[64]\ : DFN1E1C0
      port map(D => \latch_data[64]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[64]\\\);
    
    \latch_data[66]\ : DFN1E1C0
      port map(D => N_1350, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn, Q => 
        \latch_data[66]_net_1\);
    
    \Data2Fifo[30]\ : DFN1E1C0
      port map(D => \latch_data[30]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa_0, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[30]\\\);
    
    \latch4acc[10]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[10]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa_0, Q => \latch4acc[10]_net_1\);
    
    \latch_data[64]\ : DFN1E1C0
      port map(D => N_1348, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn, Q => 
        \latch_data[64]_net_1\);
    
    \latch_data[12]\ : DFN1E1C0
      port map(D => N_1602, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_3, Q
         => \latch_data[12]_net_1\);
    
    \intData2acc_RNIFHV6[4]\ : NOR3C
      port map(A => FifoRowRdOut, B => \notfirstFrame\, C => 
        \intData2acc[4]_net_1\, Y => intData2acc_RNIFHV6(4));
    
    \latch_data[48]\ : DFN1E1C0
      port map(D => N_1464, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_5, Q
         => \latch_data[48]_net_1\);
    
    \intData2acc[54]\ : DFN1E1C0
      port map(D => N_1764, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_2, Q
         => \intData2acc[54]_net_1\);
    
    \Data2Fifo[58]\ : DFN1E1C0
      port map(D => \latch_data[58]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[58]\\\);
    
    \intData2acc_RNO[36]\ : MX2
      port map(A => \latch4acc[36]_net_1\, B => 
        \intData2acc[36]_net_1\, S => N_1876, Y => N_1874);
    
    \latch_data[41]\ : DFN1E1C0
      port map(D => N_1545, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_5, Q
         => \latch_data[41]_net_1\);
    
    \intData2acc_RNITEV9[20]\ : NOR3C
      port map(A => \notfirstFrame_0\, B => 
        \intData2acc[20]_net_1\, C => FifoRowRdOut_0, Y => 
        intData2acc_RNITEV9(20));
    
    \intData2acc[0]\ : DFN1E1C0
      port map(D => N_2087, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_0, Q
         => \intData2acc[0]_net_1\);
    
    \latch_data[49]\ : DFN1E1C0
      port map(D => N_1465, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_5, Q
         => \latch_data[49]_net_1\);
    
    \intData2acc_RNO[58]\ : MX2
      port map(A => \latch4acc[58]_net_1\, B => 
        \intData2acc[58]_net_1\, S => N_1766, Y => N_1746);
    
    \intData2acc_RNIGLV6[5]\ : NOR3C
      port map(A => FifoRowRdOut, B => \notfirstFrame\, C => 
        \intData2acc[5]_net_1\, Y => intData2acc_RNIGLV6(5));
    
    \Data2Fifo[22]\ : DFN1E1C0
      port map(D => \latch_data[22]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa_0, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[22]\\\);
    
    \intData2acc_RNO[46]\ : MX2
      port map(A => \latch4acc[46]_net_1\, B => 
        \intData2acc[46]_net_1\, S => N_1876, Y => N_1821);
    
    \addSel[1]\ : DFN1C0
      port map(D => \addSel_2[1]\, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \addSel[1]_net_1\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \intData2acc[45]\ : DFN1E1C0
      port map(D => N_1820, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_2, Q
         => \intData2acc[45]_net_1\);
    
    \Data2Fifo[0]\ : DFN1E1C0
      port map(D => \latch_data[0]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa_0, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[0]\\\);
    
    \intData2acc_RNI8NV9[42]\ : NOR3C
      port map(A => FifoRowRdOut_2, B => \notfirstFrame_1\, C => 
        \intData2acc[42]_net_1\, Y => intData2acc_RNI8NV9(42));
    
    \intData2acc[36]\ : DFN1E1C0
      port map(D => N_1874, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_1, Q
         => \intData2acc[36]_net_1\);
    
    \intData2acc_RNO[25]\ : MX2
      port map(A => \latch4acc[25]_net_1\, B => 
        \intData2acc[25]_net_1\, S => N_1986, Y => N_1949);
    
    \intData2acc_RNI2KS7[28]\ : NOR3C
      port map(A => FifoRowRdOut_2, B => \notfirstFrame\, C => 
        \intData2acc[28]_net_1\, Y => intData2acc_RNI2KS7(28));
    
    \latch_data_RNO[70]\ : MX2
      port map(A => \Z\\My_adder0_3_Sum_[16]\\\, B => 
        \latch_data[70]_net_1\, S => N_15, Y => N_12);
    
    \Data2Fifo[38]\ : DFN1E1C0
      port map(D => \latch_data[38]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa_1, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[38]\\\);
    
    \latch4acc[2]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[2]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa_0, Q => \latch4acc[2]_net_1\);
    
    \latch4acc[65]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[65]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa, Q => \latch4acc[65]_net_1\);
    
    \latch4acc[18]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[18]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa_0, Q => \latch4acc[18]_net_1\);
    
    \intData2acc_RNICJ36[16]\ : NOR3C
      port map(A => FifoRowRdOut, B => \notfirstFrame\, C => 
        \intData2acc[16]_net_1\, Y => intData2acc_RNICJ36(16));
    
    \intData2acc_RNI3JV9[30]\ : NOR3C
      port map(A => FifoRowRdOut_2, B => \notfirstFrame_1\, C => 
        \intData2acc[30]_net_1\, Y => intData2acc_RNI3JV9(30));
    
    \latch_data_RNO[51]\ : MX2
      port map(A => \Z\\My_adder0_2_Sum_[15]\\\, B => 
        \latch_data[51]_net_1\, S => N_1585, Y => N_1445);
    
    \latch4acc[64]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[64]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa, Q => \latch4acc[64]_net_1\);
    
    \Data2Fifo[54]\ : DFN1E1C0
      port map(D => \latch_data[54]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[54]\\\);
    
    \Data2Fifo[67]\ : DFN1E1C0
      port map(D => \latch_data[67]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[67]\\\);
    
    \latch4acc[63]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[63]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa, Q => \latch4acc[63]_net_1\);
    
    \latch4acc[61]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[61]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa, Q => \latch4acc[61]_net_1\);
    
    \intData2acc[65]\ : DFN1E1C0
      port map(D => N_1687, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_3, Q
         => \intData2acc[65]_net_1\);
    
    \intData2acc_RNI9FV9[29]\ : NOR3C
      port map(A => FifoRowRdOut_2, B => \notfirstFrame_1\, C => 
        \intData2acc[29]_net_1\, Y => intData2acc_RNI9FV9(29));
    
    \intData2acc_RNO[31]\ : MX2
      port map(A => \latch4acc[31]_net_1\, B => 
        \intData2acc[31]_net_1\, S => N_1986, Y => N_1913);
    
    \latch_data_RNO[66]\ : MX2
      port map(A => \Z\\My_adder0_3_Sum_[12]\\\, B => 
        \latch_data[66]_net_1\, S => N_15, Y => N_1350);
    
    \latch_data_RNO[17]\ : MX2
      port map(A => \latch_data[17]_net_1\, B => 
        \Z\\My_adder0_0_Sum_[17]\\\, S => N_1657, Y => N_1562);
    
    \intData2acc_RNO[7]\ : MX2
      port map(A => \latch4acc[7]_net_1\, B => 
        \intData2acc[7]_net_1\, S => N_2090, Y => N_2055);
    
    \latch_data[33]\ : DFN1E1C0
      port map(D => N_1443, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_4, Q
         => \latch_data[33]_net_1\);
    
    \intData2acc_RNO[41]\ : MX2
      port map(A => \latch4acc[41]_net_1\, B => 
        \intData2acc[41]_net_1\, S => N_1876, Y => N_1837);
    
    \Data2Fifo[34]\ : DFN1E1C0
      port map(D => \latch_data[34]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa_1, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[34]\\\);
    
    \intData2acc_RNO[65]\ : MX2
      port map(A => \latch4acc[65]_net_1\, B => 
        \intData2acc[65]_net_1\, S => N_1766, Y => N_1687);
    
    \intData2acc_RNO[15]\ : MX2
      port map(A => \latch4acc[15]_net_1\, B => 
        \intData2acc[15]_net_1\, S => N_2090, Y => N_2003);
    
    \latch4acc[6]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[6]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa, Q => \latch4acc[6]_net_1\);
    
    \intData2acc_RNI8RV9[50]\ : NOR3C
      port map(A => FifoRowRdOut_1, B => \notfirstFrame_1\, C => 
        \intData2acc[50]_net_1\, Y => intData2acc_RNI8RV9(50));
    
    \intData2acc[24]\ : DFN1E1C0
      port map(D => N_1948, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_1, Q
         => \intData2acc[24]_net_1\);
    
    \latch_data[27]\ : DFN1E1C0
      port map(D => N_1563, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_4, Q
         => \latch_data[27]_net_1\);
    
    \latch4acc[55]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[55]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa, Q => \latch4acc[55]_net_1\);
    
    \latch_data[35]\ : DFN1E1C0
      port map(D => N_1406, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_5, Q
         => \latch_data[35]_net_1\);
    
    \latch4acc[54]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[54]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa, Q => \latch4acc[54]_net_1\);
    
    \intData2acc[4]\ : DFN1E1C0
      port map(D => N_2072, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_2, Q
         => \intData2acc[4]_net_1\);
    
    \intData2acc[42]\ : DFN1E1C0
      port map(D => N_1838, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_2, Q
         => \intData2acc[42]_net_1\);
    
    \latch_data_RNO[46]\ : MX2
      port map(A => \Z\\My_adder0_2_Sum_[10]\\\, B => 
        \latch_data[46]_net_1\, S => N_1585, Y => N_1484);
    
    \latch4acc[53]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[53]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa, Q => \latch4acc[53]_net_1\);
    
    \latch4acc[51]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[51]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa_1, Q => \latch4acc[51]_net_1\);
    
    \Data2Fifo[3]\ : DFN1E1C0
      port map(D => \latch_data[3]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa_1, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[3]\\\);
    
    \intData2acc_RNIHPV6[6]\ : NOR3C
      port map(A => FifoRowRdOut, B => \notfirstFrame\, C => 
        \intData2acc[6]_net_1\, Y => intData2acc_RNIHPV6(6));
    
    \Data2Fifo[57]\ : DFN1E1C0
      port map(D => \latch_data[57]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[57]\\\);
    
    \Data2Fifo[40]\ : DFN1E1C0
      port map(D => \latch_data[40]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa_1, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[40]\\\);
    
    \intData2acc_RNO[39]\ : MX2
      port map(A => \latch4acc[39]_net_1\, B => 
        \intData2acc[39]_net_1\, S => N_1876, Y => N_1856);
    
    \intData2acc[62]\ : DFN1E1C0
      port map(D => N_1706, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_3, Q
         => \intData2acc[62]_net_1\);
    
    \intData2acc_RNIJVV9[69]\ : NOR3C
      port map(A => FifoRowRdOut_1, B => \notfirstFrame_0\, C => 
        \intData2acc[69]_net_1\, Y => N_6);
    
    \Data2Fifo[11]\ : DFN1E1C0
      port map(D => \latch_data[11]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa_0, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[11]\\\);
    
    lvdsFifoRowRdOutEnGen : WaveGenSingleZ11
      port map(CMOS_DrvX_0_LVDSen_2 => CMOS_DrvX_0_LVDSen_2, 
        CMOS_DrvX_0_LVDSen_1 => CMOS_DrvX_0_LVDSen_1, 
        lvdsFifoRowRdOut => lvdsFifoRowRdOut, lvdsFifoRowRdOut_i
         => lvdsFifoRowRdOut_i, PLL_Test1_0_SysRst_O => 
        PLL_Test1_0_SysRst_O, PLL_Test1_0_Sys_66M_Clk => 
        PLL_Test1_0_Sys_66M_Clk);
    
    fifo_rst_n_3 : DFN1C0
      port map(D => pr_state_ns(8), CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => Main_ctl4SD_0_fifo_rst_n_3);
    
    \intData2acc_RNO[34]\ : MX2
      port map(A => \latch4acc[34]_net_1\, B => 
        \intData2acc[34]_net_1\, S => N_1986, Y => N_1895);
    
    \intData2acc_RNIARV9[54]\ : NOR3C
      port map(A => \notfirstFrame_0\, B => 
        \intData2acc[54]_net_1\, C => FifoRowRdOut_0, Y => 
        intData2acc_RNIARV9(54));
    
    \intData2acc_RNO[49]\ : MX2
      port map(A => \latch4acc[49]_net_1\, B => 
        \intData2acc[49]_net_1\, S => N_1876, Y => N_1803);
    
    \latch4acc[42]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[42]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa_1, Q => \latch4acc[42]_net_1\);
    
    \latch_data[60]\ : DFN1E1C0
      port map(D => N_1367, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn, Q => 
        \latch_data[60]_net_1\);
    
    \latch4acc[0]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[0]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa_0, Q => \latch4acc[0]_net_1\);
    
    \latch_data[17]\ : DFN1E1C0
      port map(D => N_1562, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_4, Q
         => \latch_data[17]_net_1\);
    
    \Data2Fifo[37]\ : DFN1E1C0
      port map(D => \latch_data[37]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa_1, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[37]\\\);
    
    \Data2Fifo[65]\ : DFN1E1C0
      port map(D => \latch_data[65]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[65]\\\);
    
    Data2accEnGen : WaveGenSingleZ14
      port map(PrState_2 => \PrState[4]\, PrState_0(4) => 
        \PrState_0[4]\, PLL_Test1_0_SysRst_O => 
        PLL_Test1_0_SysRst_O, PLL_Test1_0_Sys_66M_Clk => 
        PLL_Test1_0_Sys_66M_Clk, latch4acc_0_sqmuxa => 
        latch4acc_0_sqmuxa, FifoRowRdOut_1 => FifoRowRdOut_1, 
        FifoRowRdOut_0 => FifoRowRdOut_0, latch4acc_0_sqmuxa_0
         => latch4acc_0_sqmuxa_0, CMOS_DrvX_0_SDramEn_0 => 
        CMOS_DrvX_0_SDramEn_0, latch4acc_0_sqmuxa_1 => 
        latch4acc_0_sqmuxa_1);
    
    byteRdEnGen : WaveGenSingleZ8
      port map(lvdsFifoRowRdOut_i => lvdsFifoRowRdOut_i, 
        Main_ctl4SD_0_ByteRdEn => Main_ctl4SD_0_ByteRdEn, 
        PLL_Test1_0_SysRst_O => PLL_Test1_0_SysRst_O, 
        PLL_Test1_0_Sys_66M_Clk => PLL_Test1_0_Sys_66M_Clk, 
        lvdsFifoRowRdOut => lvdsFifoRowRdOut);
    
    \latch_data[42]\ : DFN1E1C0
      port map(D => N_1524, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_5, Q
         => \latch_data[42]_net_1\);
    
    \latch4acc[22]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[22]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa_0, Q => \latch4acc[22]_net_1\);
    
    \intData2acc_RNO[44]\ : MX2
      port map(A => \latch4acc[44]_net_1\, B => 
        \intData2acc[44]_net_1\, S => N_1876, Y => N_1819);
    
    \intData2acc[57]\ : DFN1E1C0
      port map(D => N_1745, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_2, Q
         => \intData2acc[57]_net_1\);
    
    \intData2acc_RNO[33]\ : MX2
      port map(A => \latch4acc[33]_net_1\, B => 
        \intData2acc[33]_net_1\, S => N_1986, Y => N_1894);
    
    \intData2acc_RNO[37]\ : MX2
      port map(A => \latch4acc[37]_net_1\, B => 
        \intData2acc[37]_net_1\, S => N_1876, Y => N_1875);
    
    \intData2acc[14]\ : DFN1E1C0
      port map(D => N_2002, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_0, Q
         => \intData2acc[14]_net_1\);
    
    \latch_data_RNO[57]\ : MX2
      port map(A => \Z\\My_adder0_3_Sum_[3]\\\, B => 
        \latch_data[57]_net_1\, S => N_15, Y => N_1387);
    
    \Data2Fifo[48]\ : DFN1E1C0
      port map(D => \latch_data[48]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa_1, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[48]\\\);
    
    \intData2acc[49]\ : DFN1E1C0
      port map(D => N_1803, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_2, Q
         => \intData2acc[49]_net_1\);
    
    \intData2acc_RNO[43]\ : MX2
      port map(A => \latch4acc[43]_net_1\, B => 
        \intData2acc[43]_net_1\, S => N_1876, Y => N_1839);
    
    \intData2acc_RNO[47]\ : MX2
      port map(A => \latch4acc[47]_net_1\, B => 
        \intData2acc[47]_net_1\, S => N_1876, Y => N_1801);
    
    \intData2acc[40]\ : DFN1E1C0
      port map(D => N_1857, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_2, Q
         => \intData2acc[40]_net_1\);
    
    \intData2acc_RNO[5]\ : MX2
      port map(A => \latch4acc[5]_net_1\, B => 
        \intData2acc[5]_net_1\, S => N_2090, Y => N_2053);
    
    \intData2acc[41]\ : DFN1E1C0
      port map(D => N_1837, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_2, Q
         => \intData2acc[41]_net_1\);
    
    \latch_data[53]\ : DFN1E1C0
      port map(D => N_1425, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_5, Q
         => \latch_data[53]_net_1\);
    
    \intData2acc_RNO[6]\ : MX2
      port map(A => \latch4acc[6]_net_1\, B => 
        \intData2acc[6]_net_1\, S => N_2090, Y => N_2054);
    
    \Data2Fifo[29]\ : DFN1E1C0
      port map(D => \latch_data[29]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa_0, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[29]\\\);
    
    \intData2acc[69]\ : DFN1E1C0
      port map(D => N_1672, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_3, Q
         => \intData2acc[69]_net_1\);
    
    \latch_data[6]\ : DFN1E1C0
      port map(D => N_1638, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn, Q => 
        \latch_data[6]_net_1\);
    
    notfirstFrame_1_sqmuxa : NOR2
      port map(A => un6_sdramenreg_net_1, B => FrameMk_0_LVDS_ok, 
        Y => \notfirstFrame_1_sqmuxa\);
    
    \latch_data[55]\ : DFN1E1C0
      port map(D => N_1408, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn, Q => 
        \latch_data[55]_net_1\);
    
    \latch_data[26]\ : DFN1E1C0
      port map(D => N_1582, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_4, Q
         => \latch_data[26]_net_1\);
    
    \intData2acc[60]\ : DFN1E1C0
      port map(D => N_1726, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_3, Q
         => \intData2acc[60]_net_1\);
    
    \Data2Fifo[44]\ : DFN1E1C0
      port map(D => \latch_data[44]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa_1, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[44]\\\);
    
    \latch_data_RNO[2]\ : MX2
      port map(A => \latch_data[2]_net_1\, B => 
        \Z\\My_adder0_0_Sum_[2]\\\, S => N_1657, Y => N_1655);
    
    \intData2acc[61]\ : DFN1E1C0
      port map(D => N_1727, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_3, Q
         => \intData2acc[61]_net_1\);
    
    \Data2Fifo[55]\ : DFN1E1C0
      port map(D => \latch_data[55]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[55]\\\);
    
    \latch_data[24]\ : DFN1E1C0
      port map(D => N_1422, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_4, Q
         => \latch_data[24]_net_1\);
    
    \latch_data_RNO[24]\ : MX2
      port map(A => \latch_data[24]_net_1\, B => 
        \Z\\My_adder0_1_Sum_[6]\\\, S => N_1546, Y => N_1422);
    
    \latch_data_RNO[13]\ : MX2
      port map(A => \latch_data[13]_net_1\, B => 
        \Z\\My_adder0_0_Sum_[13]\\\, S => N_1657, Y => N_1603);
    
    \Data2Fifo[62]\ : DFN1E1C0
      port map(D => \latch_data[62]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[62]\\\);
    
    \latch4acc[69]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[69]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa, Q => \latch4acc[69]_net_1\);
    
    \intData2acc_RNIGRV9[58]\ : NOR3C
      port map(A => FifoRowRdOut_1, B => \notfirstFrame_1\, C => 
        \intData2acc[58]_net_1\, Y => intData2acc_RNIGRV9(58));
    
    \latch_data[1]\ : DFN1E1C0
      port map(D => N_1654, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_4, Q
         => \latch_data[1]_net_1\);
    
    \latch4acc[46]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[46]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa_1, Q => \latch4acc[46]_net_1\);
    
    \intData2acc[34]\ : DFN1E1C0
      port map(D => N_1895, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_1, Q
         => \intData2acc[34]_net_1\);
    
    \intData2acc_RNO[20]\ : MX2
      port map(A => \latch4acc[20]_net_1\, B => 
        \intData2acc[20]_net_1\, S => N_1986, Y => N_1965);
    
    fifo_rst_n_6 : DFN1C0
      port map(D => pr_state_ns(8), CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => Main_ctl4SD_0_fifo_rst_n_6);
    
    \intData2acc_RNIDJ36[17]\ : NOR3C
      port map(A => FifoRowRdOut, B => \notfirstFrame\, C => 
        \intData2acc[17]_net_1\, Y => intData2acc_RNIDJ36(17));
    
    \intData2acc[27]\ : DFN1E1C0
      port map(D => N_1930, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_1, Q
         => \intData2acc[27]_net_1\);
    
    \Data2Fifo[71]\ : DFN1E1C0
      port map(D => \latch_data[71]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[71]\\\);
    
    \Data2Fifo[35]\ : DFN1E1C0
      port map(D => \latch_data[35]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa_1, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[35]\\\);
    
    \latch_data_RNO[25]\ : MX2
      port map(A => \latch_data[25]_net_1\, B => 
        \Z\\My_adder0_1_Sum_[7]\\\, S => N_1546, Y => N_1405);
    
    \latch_data[70]\ : DFN1E1C0
      port map(D => N_12, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn, Q => 
        \latch_data[70]_net_1\);
    
    \intData2acc_RNO[38]\ : MX2
      port map(A => \latch4acc[38]_net_1\, B => 
        \intData2acc[38]_net_1\, S => N_1876, Y => N_1855);
    
    \latch4acc[40]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[40]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa_1, Q => \latch4acc[40]_net_1\);
    
    \latch4acc[26]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[26]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa_0, Q => \latch4acc[26]_net_1\);
    
    \intData2acc_RNO[52]\ : MX2
      port map(A => \latch4acc[52]_net_1\, B => 
        \intData2acc[52]_net_1\, S => N_1876, Y => N_1785);
    
    \latch_data[16]\ : DFN1E1C0
      port map(D => N_1581, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_4, Q
         => \latch_data[16]_net_1\);
    
    \intData2acc[43]\ : DFN1E1C0
      port map(D => N_1839, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_2, Q
         => \intData2acc[43]_net_1\);
    
    \Data2Fifo[8]\ : DFN1E1C0
      port map(D => \latch_data[8]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[8]\\\);
    
    \intData2acc_RNIBN36[22]\ : NOR3C
      port map(A => FifoRowRdOut, B => \notfirstFrame\, C => 
        \intData2acc[22]_net_1\, Y => intData2acc_RNIBN36(22));
    
    \latch4acc[20]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[20]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa_0, Q => \latch4acc[20]_net_1\);
    
    \Data2Fifo[23]\ : DFN1E1C0
      port map(D => \latch_data[23]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa_0, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[23]\\\);
    
    \ChSel_RNO[0]\ : NOR2A
      port map(A => latch_en, B => \ChSel[0]_net_1\, Y => 
        \ChSel_3[0]\);
    
    \intData2acc_RNO[48]\ : MX2
      port map(A => \latch4acc[48]_net_1\, B => 
        \intData2acc[48]_net_1\, S => N_1876, Y => N_1802);
    
    \latch_data[14]\ : DFN1E1C0
      port map(D => N_1604, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_4, Q
         => \latch_data[14]_net_1\);
    
    \intData2acc_RNIIVV9[68]\ : NOR3C
      port map(A => FifoRowRdOut_1, B => \notfirstFrame_0\, C => 
        \intData2acc[68]_net_1\, Y => N_4);
    
    \Data2Fifo[47]\ : DFN1E1C0
      port map(D => \latch_data[47]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa_1, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[47]\\\);
    
    latchGen : WaveGenSingleZ12
      port map(PrState_4 => \PrState[4]\, PrState_0(4) => 
        \PrState_0[4]\, latch_en => latch_en, FifoRowRdOut => 
        FifoRowRdOut, FifoRowRdOut_0 => FifoRowRdOut_0, 
        PLL_Test1_0_SysRst_O => PLL_Test1_0_SysRst_O, 
        FifoRowRdOut_i => FifoRowRdOut_i, PLL_Test1_0_Sys_66M_Clk
         => PLL_Test1_0_Sys_66M_Clk);
    
    \latch4acc[59]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[59]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa, Q => \latch4acc[59]_net_1\);
    
    \latch4acc[35]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[35]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa_1, Q => \latch4acc[35]_net_1\);
    
    \latch4acc[34]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[34]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa_1, Q => \latch4acc[34]_net_1\);
    
    \intData2acc_RNO[3]\ : MX2
      port map(A => \latch4acc[3]_net_1\, B => 
        \intData2acc[3]_net_1\, S => N_2090, Y => N_2071);
    
    \latch4acc[3]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[3]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa_1, Q => \latch4acc[3]_net_1\);
    
    \latch4acc[33]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[33]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa_1, Q => \latch4acc[33]_net_1\);
    
    \latch4acc[31]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[31]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa_1, Q => \latch4acc[31]_net_1\);
    
    \Data2Fifo[52]\ : DFN1E1C0
      port map(D => \latch_data[52]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa_1, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[52]\\\);
    
    \ChSel_RNITABA[1]\ : OR2B
      port map(A => \ChSel[1]_net_1\, B => \ChSel[0]_net_1\, Y
         => N_15);
    
    \intData2acc[63]\ : DFN1E1C0
      port map(D => N_1707, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_3, Q
         => \intData2acc[63]_net_1\);
    
    \intData2acc_RNO[60]\ : MX2
      port map(A => \latch4acc[60]_net_1\, B => 
        \intData2acc[60]_net_1\, S => N_1766, Y => N_1726);
    
    \intData2acc_RNO[10]\ : MX2
      port map(A => \latch4acc[10]_net_1\, B => 
        \intData2acc[10]_net_1\, S => N_2090, Y => N_2038);
    
    fifo_rdGen : WaveGenSingleZ16
      port map(PrState_2 => \PrState[4]\, PrState_0(4) => 
        \PrState_0[4]\, PLL_Test1_0_SysRst_O => 
        PLL_Test1_0_SysRst_O, PLL_Test1_0_Sys_66M_Clk => 
        PLL_Test1_0_Sys_66M_Clk, lvds_fifoRd => lvds_fifoRd, 
        Main_ctl4SD_0_fifo_rd => Main_ctl4SD_0_fifo_rd, 
        FifoRowRdOut_1 => FifoRowRdOut_1, FifoRowRdOut_0 => 
        FifoRowRdOut_0);
    
    \latch_data_RNO[10]\ : MX2
      port map(A => \latch_data[10]_net_1\, B => 
        \Z\\My_adder0_0_Sum_[10]\\\, S => N_1657, Y => N_1621);
    
    \latch_data_RNO[29]\ : MX2
      port map(A => \latch_data[29]_net_1\, B => 
        \Z\\My_adder0_1_Sum_[11]\\\, S => N_1546, Y => N_1523);
    
    \intData2acc_RNO[26]\ : MX2
      port map(A => \latch4acc[26]_net_1\, B => 
        \intData2acc[26]_net_1\, S => N_1986, Y => N_1929);
    
    \intData2acc[48]\ : DFN1E1C0
      port map(D => N_1802, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_2, Q
         => \intData2acc[48]_net_1\);
    
    \latch_data_RNO[18]\ : MX2
      port map(A => \latch_data[18]_net_1\, B => 
        \Z\\My_adder0_1_Sum_[0]\\\, S => N_1546, Y => N_1542);
    
    \latch_data[47]\ : DFN1E1C0
      port map(D => N_1485, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_5, Q
         => \latch_data[47]_net_1\);
    
    \latch4acc[48]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[48]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa_1, Q => \latch4acc[48]_net_1\);
    
    \latch_data[38]\ : DFN1E1C0
      port map(D => N_1564, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_5, Q
         => \latch_data[38]_net_1\);
    
    \ChSel[1]\ : DFN1C0
      port map(D => \ChSel_3[1]\, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \ChSel[1]_net_1\);
    
    \latch_data_RNO[53]\ : MX2
      port map(A => \Z\\My_adder0_2_Sum_[17]\\\, B => 
        \latch_data[53]_net_1\, S => N_1585, Y => N_1425);
    
    \latch_data_RNO[12]\ : MX2
      port map(A => \latch_data[12]_net_1\, B => 
        \Z\\My_adder0_0_Sum_[12]\\\, S => N_1657, Y => N_1602);
    
    \latch_data[31]\ : DFN1E1C0
      port map(D => N_1483, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_4, Q
         => \latch_data[31]_net_1\);
    
    \intData2acc[17]\ : DFN1E1C0
      port map(D => N_1983, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_1, Q
         => \intData2acc[17]_net_1\);
    
    \latch4acc[28]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[28]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa_0, Q => \latch4acc[28]_net_1\);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    \latch_data[39]\ : DFN1E1C0
      port map(D => N_1565, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_5, Q
         => \latch_data[39]_net_1\);
    
    \Data2Fifo[26]\ : DFN1E1C0
      port map(D => \latch_data[26]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa_0, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[26]\\\);
    
    \Data2Fifo[32]\ : DFN1E1C0
      port map(D => \latch_data[32]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa_1, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[32]\\\);
    
    \latch_data_RNO[34]\ : MX2
      port map(A => \latch_data[34]_net_1\, B => 
        \Z\\My_adder0_1_Sum_[16]\\\, S => N_1546, Y => N_1423);
    
    \intData2acc[68]\ : DFN1E1C0
      port map(D => N_1671, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_3, Q
         => \intData2acc[68]_net_1\);
    
    FifoRowRdOutGen : WaveGenSingleZ17
      port map(FifoRowRdOut => FifoRowRdOut, 
        CMOS_DrvX_0_SDramEn_0 => CMOS_DrvX_0_SDramEn_0, 
        FifoRowRdOut_i => FifoRowRdOut_i, FifoRowRdOut_0 => 
        FifoRowRdOut_0, FifoRowRdOut_1 => FifoRowRdOut_1, 
        PLL_Test1_0_SysRst_O => PLL_Test1_0_SysRst_O, 
        PLL_Test1_0_Sys_66M_Clk => PLL_Test1_0_Sys_66M_Clk, 
        FifoRowRdOut_2 => FifoRowRdOut_2);
    
    \intData2acc_RNIFVV9[65]\ : NOR3C
      port map(A => FifoRowRdOut_1, B => \notfirstFrame_0\, C => 
        \intData2acc[65]_net_1\, Y => intData2acc_RNIFVV9(65));
    
    \latch4acc[70]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[70]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa, Q => \latch4acc[70]_net_1\);
    
    \intData2acc_RNO[66]\ : MX2
      port map(A => \latch4acc[66]_net_1\, B => 
        \intData2acc[66]_net_1\, S => N_1766, Y => N_1688);
    
    \intData2acc_RNO[16]\ : MX2
      port map(A => \latch4acc[16]_net_1\, B => 
        \intData2acc[16]_net_1\, S => N_2090, Y => N_2004);
    
    \intData2acc_RNIDRV9[56]\ : NOR3C
      port map(A => FifoRowRdOut_1, B => \notfirstFrame_0\, C => 
        \intData2acc[56]_net_1\, Y => intData2acc_RNIDRV9(56));
    
    \latch4acc[67]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[67]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa, Q => \latch4acc[67]_net_1\);
    
    fifo_rst_n_1 : DFN1C0
      port map(D => pr_state_ns(8), CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => Main_ctl4SD_0_fifo_rst_n_1);
    
    \latch_data_RNO[35]\ : MX2
      port map(A => \latch_data[35]_net_1\, B => 
        \Z\\My_adder0_1_Sum_[17]\\\, S => N_1546, Y => N_1406);
    
    \latch_data[63]\ : DFN1E1C0
      port map(D => N_1370, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn, Q => 
        \latch_data[63]_net_1\);
    
    \latch4acc[8]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[8]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa, Q => \latch4acc[8]_net_1\);
    
    \intData2acc_RNO[21]\ : MX2
      port map(A => \latch4acc[21]_net_1\, B => 
        \intData2acc[21]_net_1\, S => N_1986, Y => N_1966);
    
    \Data2Fifo[10]\ : DFN1E1C0
      port map(D => \latch_data[10]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa_0, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[10]\\\);
    
    \Data2Fifo[1]\ : DFN1E1C0
      port map(D => \latch_data[1]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa_0, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[1]\\\);
    
    \latch_data[20]\ : DFN1E1C0
      port map(D => N_1502, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_4, Q
         => \latch_data[20]_net_1\);
    
    \addSel_RNILVIF_2[1]\ : OR2
      port map(A => \addSel[1]_net_1\, B => \addSel[0]_net_1\, Y
         => N_2090);
    
    \intData2acc_RNI7JV9[37]\ : NOR3C
      port map(A => \notfirstFrame_0\, B => 
        \intData2acc[37]_net_1\, C => FifoRowRdOut_0, Y => 
        intData2acc_RNI7JV9_3);
    
    \Data2Fifo[45]\ : DFN1E1C0
      port map(D => \latch_data[45]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa_1, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[45]\\\);
    
    \latch_data[65]\ : DFN1E1C0
      port map(D => N_1349, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn, Q => 
        \latch_data[65]_net_1\);
    
    \intData2acc_RNO[0]\ : MX2
      port map(A => \latch4acc[0]_net_1\, B => 
        \intData2acc[0]_net_1\, S => N_2090, Y => N_2087);
    
    \latch_data_RNO[21]\ : MX2
      port map(A => \latch_data[21]_net_1\, B => 
        \Z\\My_adder0_1_Sum_[3]\\\, S => N_1546, Y => N_1482);
    
    \intData2acc_RNIK507[9]\ : NOR3C
      port map(A => FifoRowRdOut, B => \notfirstFrame\, C => 
        \intData2acc[9]_net_1\, Y => intData2acc_RNIK507(9));
    
    \intData2acc_RNIENV9[48]\ : NOR3C
      port map(A => FifoRowRdOut_2, B => \notfirstFrame_1\, C => 
        \intData2acc[48]_net_1\, Y => intData2acc_RNIENV9(48));
    
    \latch_data_RNO[50]\ : MX2
      port map(A => \Z\\My_adder0_2_Sum_[14]\\\, B => 
        \latch_data[50]_net_1\, S => N_1585, Y => N_1444);
    
    \latch_data_RNO[58]\ : MX2
      port map(A => \Z\\My_adder0_3_Sum_[4]\\\, B => 
        \latch_data[58]_net_1\, S => N_15, Y => N_1388);
    
    \intData2acc_RNIGRV9[59]\ : NOR3C
      port map(A => FifoRowRdOut_1, B => \notfirstFrame_0\, C => 
        \intData2acc[59]_net_1\, Y => intData2acc_RNIGRV9(59));
    
    \intData2acc[37]\ : DFN1E1C0
      port map(D => N_1875, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_2, Q
         => \intData2acc[37]_net_1\);
    
    \latch_data[4]\ : DFN1E1C0
      port map(D => N_1636, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_5, Q
         => \latch_data[4]_net_1\);
    
    \Data2Fifo[7]\ : DFN1E1C0
      port map(D => \latch_data[7]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[7]\\\);
    
    \Data2Fifo[69]\ : DFN1E1C0
      port map(D => \latch_data[69]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[69]\\\);
    
    \latch_data_RNO[52]\ : MX2
      port map(A => \Z\\My_adder0_2_Sum_[16]\\\, B => 
        \latch_data[52]_net_1\, S => N_1585, Y => N_1424);
    
    \addSel_RNO[1]\ : XA1B
      port map(A => \addSel[0]_net_1\, B => \addSel[1]_net_1\, C
         => CMOS_DrvX_0_AdcEn, Y => \addSel_2[1]\);
    
    \latch_data_RNO[39]\ : MX2
      port map(A => \Z\\My_adder0_2_Sum_[3]\\\, B => 
        \latch_data[39]_net_1\, S => N_1585, Y => N_1565);
    
    \latch4acc[57]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[57]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa, Q => \latch4acc[57]_net_1\);
    
    \latch4acc[15]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[15]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa_0, Q => \latch4acc[15]_net_1\);
    
    \intData2acc_RNO[61]\ : MX2
      port map(A => \latch4acc[61]_net_1\, B => 
        \intData2acc[61]_net_1\, S => N_1766, Y => N_1727);
    
    \intData2acc_RNO[11]\ : MX2
      port map(A => \latch4acc[11]_net_1\, B => 
        \intData2acc[11]_net_1\, S => N_2090, Y => N_2019);
    
    \Data2Fifo[18]\ : DFN1E1C0
      port map(D => \latch_data[18]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa_0, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[18]\\\);
    
    \latch4acc[14]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[14]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa_0, Q => \latch4acc[14]_net_1\);
    
    \intData2acc[46]\ : DFN1E1C0
      port map(D => N_1821, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_2, Q
         => \intData2acc[46]_net_1\);
    
    \latch_data[58]\ : DFN1E1C0
      port map(D => N_1388, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn, Q => 
        \latch_data[58]_net_1\);
    
    \latch_data[46]\ : DFN1E1C0
      port map(D => N_1484, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_5, Q
         => \latch_data[46]_net_1\);
    
    \latch4acc[13]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[13]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa_0, Q => \latch4acc[13]_net_1\);
    
    \latch4acc[11]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[11]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa_0, Q => \latch4acc[11]_net_1\);
    
    \intData2acc_RNO[29]\ : MX2
      port map(A => \latch4acc[29]_net_1\, B => 
        \intData2acc[29]_net_1\, S => N_1986, Y => N_1911);
    
    \ChSel_RNO[1]\ : XA1
      port map(A => \ChSel[0]_net_1\, B => \ChSel[1]_net_1\, C
         => latch_en, Y => \ChSel_3[1]\);
    
    \latch_data[10]\ : DFN1E1C0
      port map(D => N_1621, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_3, Q
         => \latch_data[10]_net_1\);
    
    \intData2acc_RNO[70]\ : MX2
      port map(A => \latch4acc[70]_net_1\, B => 
        \intData2acc[70]_net_1\, S => N_1766, Y => N_1673);
    
    \intData2acc[55]\ : DFN1E1C0
      port map(D => N_1765, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_2, Q
         => \intData2acc[55]_net_1\);
    
    \latch_data[51]\ : DFN1E1C0
      port map(D => N_1445, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_5, Q
         => \latch_data[51]_net_1\);
    
    lvds_fifoRdGen : WaveGenSingleZ10
      port map(lvds_fifoRd => lvds_fifoRd, PLL_Test1_0_SysRst_O
         => PLL_Test1_0_SysRst_O, PLL_Test1_0_Sys_66M_Clk => 
        PLL_Test1_0_Sys_66M_Clk, lvdsFifoRowRdOut => 
        lvdsFifoRowRdOut);
    
    \latch_data[59]\ : DFN1E1C0
      port map(D => N_1389, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn, Q => 
        \latch_data[59]_net_1\);
    
    \latch_data[44]\ : DFN1E1C0
      port map(D => N_1504, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_5, Q
         => \latch_data[44]_net_1\);
    
    fifo_wrGen : WaveGenSingleZ15
      port map(Main_ctl4SD_0_Fifo_wr => Main_ctl4SD_0_Fifo_wr, 
        PLL_Test1_0_SysRst_O => PLL_Test1_0_SysRst_O, 
        PLL_Test1_0_Sys_66M_Clk => PLL_Test1_0_Sys_66M_Clk, 
        FifoRowRdOut_1 => FifoRowRdOut_1, FifoRowRdOut_0 => 
        FifoRowRdOut_0);
    
    \latch_data_RNO[16]\ : MX2
      port map(A => \latch_data[16]_net_1\, B => 
        \Z\\My_adder0_0_Sum_[16]\\\, S => N_1657, Y => N_1581);
    
    \intData2acc_RNO[24]\ : MX2
      port map(A => \latch4acc[24]_net_1\, B => 
        \intData2acc[24]_net_1\, S => N_1986, Y => N_1948);
    
    \intData2acc[66]\ : DFN1E1C0
      port map(D => N_1688, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_3, Q
         => \intData2acc[66]_net_1\);
    
    \latch_data_RNO[64]\ : MX2
      port map(A => \Z\\My_adder0_3_Sum_[10]\\\, B => 
        \latch_data[64]_net_1\, S => N_15, Y => N_1348);
    
    \latch4acc[1]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[1]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa_0, Q => \latch4acc[1]_net_1\);
    
    \Data2Fifo[42]\ : DFN1E1C0
      port map(D => \latch_data[42]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa_1, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[42]\\\);
    
    \intData2acc_RNO[23]\ : MX2
      port map(A => \latch4acc[23]_net_1\, B => 
        \intData2acc[23]_net_1\, S => N_1986, Y => N_1947);
    
    \Data2Fifo[14]\ : DFN1E1C0
      port map(D => \latch_data[14]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa_0, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[14]\\\);
    
    \intData2acc_RNO[27]\ : MX2
      port map(A => \latch4acc[27]_net_1\, B => 
        \intData2acc[27]_net_1\, S => N_1986, Y => N_1930);
    
    \intData2acc_RNI2BV9[18]\ : NOR3C
      port map(A => \notfirstFrame_0\, B => 
        \intData2acc[18]_net_1\, C => FifoRowRdOut_0, Y => 
        intData2acc_RNI2BV9(18));
    
    \latch_data[32]\ : DFN1E1C0
      port map(D => N_1463, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_4, Q
         => \latch_data[32]_net_1\);
    
    \latch_data_RNO[4]\ : MX2
      port map(A => \latch_data[4]_net_1\, B => 
        \Z\\My_adder0_0_Sum_[4]\\\, S => N_1657, Y => N_1636);
    
    \Data2Fifo[59]\ : DFN1E1C0
      port map(D => \latch_data[59]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[59]\\\);
    
    \latch4acc[39]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[39]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa_1, Q => \latch4acc[39]_net_1\);
    
    \intData2acc_RNO[69]\ : MX2
      port map(A => \latch4acc[69]_net_1\, B => 
        \intData2acc[69]_net_1\, S => N_1766, Y => N_1672);
    
    \intData2acc_RNO[19]\ : MX2
      port map(A => \latch4acc[19]_net_1\, B => 
        \intData2acc[19]_net_1\, S => N_1986, Y => N_1985);
    
    fifo_rst_n_5 : DFN1C0
      port map(D => pr_state_ns(8), CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => Main_ctl4SD_0_fifo_rst_n_5);
    
    \Data2Fifo[2]\ : DFN1E1C0
      port map(D => \latch_data[2]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa_0, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[2]\\\);
    
    \Data2Fifo[21]\ : DFN1E1C0
      port map(D => \latch_data[21]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa_0, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[21]\\\);
    
    \latch_data_RNO[65]\ : MX2
      port map(A => \Z\\My_adder0_3_Sum_[11]\\\, B => 
        \latch_data[65]_net_1\, S => N_15, Y => N_1349);
    
    \Data2Fifo[63]\ : DFN1E1C0
      port map(D => \latch_data[63]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[63]\\\);
    
    Data2fifoENGen : WaveGenSingleZ13
      port map(PLL_Test1_0_SysRst_O => PLL_Test1_0_SysRst_O, 
        PLL_Test1_0_Sys_66M_Clk => PLL_Test1_0_Sys_66M_Clk, 
        FifoRowRdOut => FifoRowRdOut, Data2Fifo_0_sqmuxa => 
        Data2Fifo_0_sqmuxa, FifoRowRdOut_1 => FifoRowRdOut_1, 
        FifoRowRdOut_0 => FifoRowRdOut_0, Data2Fifo_0_sqmuxa_0
         => Data2Fifo_0_sqmuxa_0, CMOS_DrvX_0_SDramEn_0 => 
        CMOS_DrvX_0_SDramEn_0, Data2Fifo_0_sqmuxa_1 => 
        Data2Fifo_0_sqmuxa_1);
    
    \latch_data_RNO[44]\ : MX2
      port map(A => \Z\\My_adder0_2_Sum_[8]\\\, B => 
        \latch_data[44]_net_1\, S => N_1585, Y => N_1504);
    
    \intData2acc_RNI8JV9[35]\ : NOR3C
      port map(A => FifoRowRdOut_2, B => \notfirstFrame_1\, C => 
        \intData2acc[35]_net_1\, Y => intData2acc_RNI8JV9(35));
    
    \Data2Fifo[70]\ : DFN1E1C0
      port map(D => \latch_data[70]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[70]\\\);
    
    \intData2acc_RNO[64]\ : MX2
      port map(A => \latch4acc[64]_net_1\, B => 
        \intData2acc[64]_net_1\, S => N_1766, Y => N_1708);
    
    \intData2acc_RNO[14]\ : MX2
      port map(A => \latch4acc[14]_net_1\, B => 
        \intData2acc[14]_net_1\, S => N_2090, Y => N_2002);
    
    \intData2acc_RNI6NV9[40]\ : NOR3C
      port map(A => FifoRowRdOut_2, B => \notfirstFrame_1\, C => 
        \intData2acc[40]_net_1\, Y => intData2acc_RNI6NV9(40));
    
    \ChSel_RNITABA_0[1]\ : OR2A
      port map(A => \ChSel[1]_net_1\, B => \ChSel[0]_net_1\, Y
         => N_1585);
    
    \latch_data_RNO[31]\ : MX2
      port map(A => \latch_data[31]_net_1\, B => 
        \Z\\My_adder0_1_Sum_[13]\\\, S => N_1546, Y => N_1483);
    
    \intData2acc[52]\ : DFN1E1C0
      port map(D => N_1785, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_2, Q
         => \intData2acc[52]_net_1\);
    
    \intData2acc_RNO[32]\ : MX2
      port map(A => \latch4acc[32]_net_1\, B => 
        \intData2acc[32]_net_1\, S => N_1986, Y => N_1893);
    
    \intData2acc_RNIDVV9[63]\ : NOR3C
      port map(A => FifoRowRdOut_1, B => \notfirstFrame_0\, C => 
        \intData2acc[63]_net_1\, Y => intData2acc_RNIDVV9(63));
    
    \intData2acc_RNIJ107[8]\ : NOR3C
      port map(A => FifoRowRdOut, B => \notfirstFrame\, C => 
        \intData2acc[8]_net_1\, Y => intData2acc_RNIJ107(8));
    
    \Data2Fifo[39]\ : DFN1E1C0
      port map(D => \latch_data[39]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa_1, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[39]\\\);
    
    \latch_data_RNO[27]\ : MX2
      port map(A => \latch_data[27]_net_1\, B => 
        \Z\\My_adder0_1_Sum_[9]\\\, S => N_1546, Y => N_1563);
    
    \intData2acc_RNO[63]\ : MX2
      port map(A => \latch4acc[63]_net_1\, B => 
        \intData2acc[63]_net_1\, S => N_1766, Y => N_1707);
    
    \intData2acc_RNO[13]\ : MX2
      port map(A => \latch4acc[13]_net_1\, B => 
        \intData2acc[13]_net_1\, S => N_2090, Y => N_2021);
    
    \intData2acc[2]\ : DFN1E1C0
      port map(D => N_2070, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_1, Q
         => \intData2acc[2]_net_1\);
    
    \intData2acc_RNO[67]\ : MX2
      port map(A => \latch4acc[67]_net_1\, B => 
        \intData2acc[67]_net_1\, S => N_1766, Y => N_1689);
    
    \intData2acc_RNO[17]\ : MX2
      port map(A => \latch4acc[17]_net_1\, B => 
        \intData2acc[17]_net_1\, S => N_2090, Y => N_1983);
    
    \latch_data_RNO[45]\ : MX2
      port map(A => \Z\\My_adder0_2_Sum_[9]\\\, B => 
        \latch_data[45]_net_1\, S => N_1585, Y => N_1505);
    
    \intData2acc[9]\ : DFN1E1C0
      port map(D => N_2037, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_3, Q
         => \intData2acc[9]_net_1\);
    
    \intData2acc_RNO[42]\ : MX2
      port map(A => \latch4acc[42]_net_1\, B => 
        \intData2acc[42]_net_1\, S => N_1876, Y => N_1838);
    
    \intData2acc[25]\ : DFN1E1C0
      port map(D => N_1949, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_1, Q
         => \intData2acc[25]_net_1\);
    
    \intData2acc_RNO[55]\ : MX2
      port map(A => \latch4acc[55]_net_1\, B => 
        \intData2acc[55]_net_1\, S => N_1766, Y => N_1765);
    
    \Data2Fifo[17]\ : DFN1E1C0
      port map(D => \latch_data[17]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa_0, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[17]\\\);
    
    \latch_data_RNO[56]\ : MX2
      port map(A => \Z\\My_adder0_3_Sum_[2]\\\, B => 
        \latch_data[56]_net_1\, S => N_15, Y => N_1386);
    
    \latch_data_RNO[69]\ : MX2
      port map(A => \Z\\My_adder0_3_Sum_[15]\\\, B => 
        \latch_data[69]_net_1\, S => N_15, Y => N_10);
    
    \Data2Fifo[66]\ : DFN1E1C0
      port map(D => \latch_data[66]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[66]\\\);
    
    \latch4acc[62]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[62]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa, Q => \latch4acc[62]_net_1\);
    
    \intData2acc_RNI1KS7[27]\ : NOR3C
      port map(A => FifoRowRdOut_2, B => \notfirstFrame\, C => 
        \intData2acc[27]_net_1\, Y => intData2acc_RNI1KS7(27));
    
    \intData2acc_RNO[71]\ : MX2
      port map(A => \latch4acc[71]_net_1\, B => 
        \intData2acc[71]_net_1\, S => N_1766, Y => N_2089);
    
    \Data2Fifo[53]\ : DFN1E1C0
      port map(D => \latch_data[53]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[53]\\\);
    
    \latch4acc[4]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[4]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa_1, Q => \latch4acc[4]_net_1\);
    
    \latch4acc[9]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[9]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa, Q => \latch4acc[9]_net_1\);
    
    \intData2acc_RNO[28]\ : MX2
      port map(A => \latch4acc[28]_net_1\, B => 
        \intData2acc[28]_net_1\, S => N_1986, Y => N_1931);
    
    \intData2acc[70]\ : DFN1E1C0
      port map(D => N_1673, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_3, Q
         => \intData2acc[70]_net_1\);
    
    \latch_data_RNO[49]\ : MX2
      port map(A => \Z\\My_adder0_2_Sum_[13]\\\, B => 
        \latch_data[49]_net_1\, S => N_1585, Y => N_1465);
    
    \intData2acc_RNICJV9[39]\ : NOR3C
      port map(A => FifoRowRdOut_2, B => \notfirstFrame_1\, C => 
        \intData2acc[39]_net_1\, Y => intData2acc_RNICJV9(39));
    
    \intData2acc_RNI11RA[2]\ : NOR3C
      port map(A => \notfirstFrame_0\, B => 
        \intData2acc[2]_net_1\, C => FifoRowRdOut_0, Y => 
        intData2acc_RNI11RA(2));
    
    \intData2acc[71]\ : DFN1E1C0
      port map(D => N_2089, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_3, Q
         => \intData2acc[71]_net_1\);
    
    \intData2acc[59]\ : DFN1E1C0
      port map(D => N_1725, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_3, Q
         => \intData2acc[59]_net_1\);
    
    \intData2acc_RNIERV9[57]\ : NOR3C
      port map(A => FifoRowRdOut_1, B => \notfirstFrame_0\, C => 
        \intData2acc[57]_net_1\, Y => intData2acc_RNIERV9(57));
    
    \latch_data[52]\ : DFN1E1C0
      port map(D => N_1424, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_5, Q
         => \latch_data[52]_net_1\);
    
    \intData2acc_RNI8J36[12]\ : NOR3C
      port map(A => FifoRowRdOut, B => \notfirstFrame\, C => 
        \intData2acc[12]_net_1\, Y => intData2acc_RNI8J36(12));
    
    \intData2acc_RNIEDV6[3]\ : NOR3C
      port map(A => FifoRowRdOut, B => \notfirstFrame\, C => 
        \intData2acc[3]_net_1\, Y => intData2acc_RNIEDV6(3));
    
    \intData2acc[7]\ : DFN1E1C0
      port map(D => N_2055, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_3, Q
         => \intData2acc[7]_net_1\);
    
    \intData2acc[50]\ : DFN1E1C0
      port map(D => N_1783, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_2, Q
         => \intData2acc[50]_net_1\);
    
    \Data2Fifo[33]\ : DFN1E1C0
      port map(D => \latch_data[33]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa_1, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[33]\\\);
    
    \latch_data[40]\ : DFN1E1C0
      port map(D => N_1544, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_5, Q
         => \latch_data[40]_net_1\);
    
    \intData2acc[51]\ : DFN1E1C0
      port map(D => N_1784, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_2, Q
         => \intData2acc[51]_net_1\);
    
    \latch_data[23]\ : DFN1E1C0
      port map(D => N_1442, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_4, Q
         => \latch_data[23]_net_1\);
    
    \latch_data[0]\ : DFN1E1C0
      port map(D => N_1653, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_3, Q
         => \latch_data[0]_net_1\);
    
    \intData2acc[15]\ : DFN1E1C0
      port map(D => N_2003, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_0, Q
         => \intData2acc[15]_net_1\);
    
    \latch4acc[52]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[52]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa_1, Q => \latch4acc[52]_net_1\);
    
    \intData2acc_RNIBVV9[61]\ : NOR3C
      port map(A => FifoRowRdOut_1, B => \notfirstFrame_0\, C => 
        \intData2acc[61]_net_1\, Y => intData2acc_RNIBVV9(61));
    
    \intData2acc[22]\ : DFN1E1C0
      port map(D => N_1967, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_1, Q
         => \intData2acc[22]_net_1\);
    
    \addSel_RNILVIF_1[1]\ : OR2A
      port map(A => \addSel[0]_net_1\, B => \addSel[1]_net_1\, Y
         => N_1986);
    
    \latch_data[68]\ : DFN1E1C0
      port map(D => N_8, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn, Q => 
        \latch_data[68]_net_1\);
    
    \intData2acc_RNO[8]\ : MX2
      port map(A => \latch4acc[8]_net_1\, B => 
        \intData2acc[8]_net_1\, S => N_2090, Y => N_2036);
    
    \latch_data[5]\ : DFN1E1C0
      port map(D => N_1637, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn, Q => 
        \latch_data[5]_net_1\);
    
    \Data2Fifo[56]\ : DFN1E1C0
      port map(D => \latch_data[56]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[56]\\\);
    
    \latch4acc[37]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[37]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa_1, Q => \latch4acc[37]_net_1\);
    
    \latch_data[61]\ : DFN1E1C0
      port map(D => N_1368, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn, Q => 
        \latch_data[61]_net_1\);
    
    \latch4acc[19]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[19]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa_0, Q => \latch4acc[19]_net_1\);
    
    \intData2acc_RNO[68]\ : MX2
      port map(A => \latch4acc[68]_net_1\, B => 
        \intData2acc[68]_net_1\, S => N_1766, Y => N_1671);
    
    \intData2acc_RNO[18]\ : MX2
      port map(A => \latch4acc[18]_net_1\, B => 
        \intData2acc[18]_net_1\, S => N_1986, Y => N_1984);
    
    \Data2Fifo[9]\ : DFN1E1C0
      port map(D => \latch_data[9]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[9]\\\);
    
    \latch_data[69]\ : DFN1E1C0
      port map(D => N_10, CLK => PLL_Test1_0_Sys_66M_Clk, CLR => 
        PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn, Q => 
        \latch_data[69]_net_1\);
    
    \latch_data[25]\ : DFN1E1C0
      port map(D => N_1405, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_4, Q
         => \latch_data[25]_net_1\);
    
    \latch_data_RNO[61]\ : MX2
      port map(A => \Z\\My_adder0_3_Sum_[7]\\\, B => 
        \latch_data[61]_net_1\, S => N_15, Y => N_1368);
    
    \latch_data_RNO[37]\ : MX2
      port map(A => \Z\\My_adder0_2_Sum_[1]\\\, B => 
        \latch_data[37]_net_1\, S => N_1585, Y => N_1584);
    
    \addSel_RNILVIF_0[1]\ : OR2A
      port map(A => \addSel[1]_net_1\, B => \addSel[0]_net_1\, Y
         => N_1876);
    
    \latch_data[37]\ : DFN1E1C0
      port map(D => N_1584, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_5, Q
         => \latch_data[37]_net_1\);
    
    \intData2acc_RNIAJ36[14]\ : NOR3C
      port map(A => FifoRowRdOut, B => \notfirstFrame\, C => 
        \intData2acc[14]_net_1\, Y => intData2acc_RNIAJ36(14));
    
    \intData2acc_RNI6JV9[36]\ : NOR3C
      port map(A => \notfirstFrame_0\, B => 
        \intData2acc[36]_net_1\, C => FifoRowRdOut_0, Y => 
        intData2acc_RNI6JV9_3);
    
    \Data2Fifo[15]\ : DFN1E1C0
      port map(D => \latch_data[15]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa_0, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[15]\\\);
    
    \intData2acc[44]\ : DFN1E1C0
      port map(D => N_1819, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_2, Q
         => \intData2acc[44]_net_1\);
    
    \Data2Fifo[49]\ : DFN1E1C0
      port map(D => \latch_data[49]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa_1, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[49]\\\);
    
    \Data2Fifo[36]\ : DFN1E1C0
      port map(D => \latch_data[36]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => Data2Fifo_0_sqmuxa_1, Q => 
        \Z\\Main_ctl4SD_0_Data2Fifo_[36]\\\);
    
    \latch4acc[66]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[66]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa, Q => \latch4acc[66]_net_1\);
    
    \intData2acc_RNI0TQA[1]\ : NOR3C
      port map(A => \notfirstFrame_0\, B => 
        \intData2acc[1]_net_1\, C => FifoRowRdOut_0, Y => 
        intData2acc_RNI0TQA(1));
    
    \latch_data[13]\ : DFN1E1C0
      port map(D => N_1603, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_4, Q
         => \latch_data[13]_net_1\);
    
    \intData2acc_RNI6JV9[33]\ : NOR3C
      port map(A => FifoRowRdOut_2, B => \notfirstFrame_1\, C => 
        \intData2acc[33]_net_1\, Y => intData2acc_RNI6JV9_0);
    
    \latch_data_RNO[41]\ : MX2
      port map(A => \Z\\My_adder0_2_Sum_[5]\\\, B => 
        \latch_data[41]_net_1\, S => N_1585, Y => N_1545);
    
    \latch_data[7]\ : DFN1E1C0
      port map(D => N_1639, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn, Q => 
        \latch_data[7]_net_1\);
    
    \latch4acc[60]\ : DFN1E1C0
      port map(D => \Z\\Fifo_rd_0_Q_[60]\\\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => latch4acc_0_sqmuxa, Q => \latch4acc[60]_net_1\);
    
    \intData2acc_RNIAVV9[60]\ : NOR3C
      port map(A => FifoRowRdOut_1, B => \notfirstFrame_0\, C => 
        \intData2acc[60]_net_1\, Y => intData2acc_RNIAVV9(60));
    
    \latch_data[2]\ : DFN1E1C0
      port map(D => N_1655, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_4, Q
         => \latch_data[2]_net_1\);
    
    \latch_data[15]\ : DFN1E1C0
      port map(D => N_1605, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_4, Q
         => \latch_data[15]_net_1\);
    
    \intData2acc[64]\ : DFN1E1C0
      port map(D => N_1708, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_3, Q
         => \intData2acc[64]_net_1\);
    
    \intData2acc[12]\ : DFN1E1C0
      port map(D => N_2020, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_0, Q
         => \intData2acc[12]_net_1\);
    
    \latch_data_RNO[23]\ : MX2
      port map(A => \latch_data[23]_net_1\, B => 
        \Z\\My_adder0_1_Sum_[5]\\\, S => N_1546, Y => N_1442);
    
    \intData2acc[29]\ : DFN1E1C0
      port map(D => N_1911, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_1, Q
         => \intData2acc[29]_net_1\);
    
    \intData2acc[53]\ : DFN1E1C0
      port map(D => N_1763, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => CMOS_DrvX_0_SDramEn_2, Q
         => \intData2acc[53]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3;
use proasic3.all;

entity Fifo_rd_1 is

    port( \Z\\Fifo_rd_0_Q_[27]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[23]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[69]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[1]\\\               : out   std_logic;
          \Z\\Fifo_rd_0_Q_[67]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[4]\\\               : out   std_logic;
          \Z\\Fifo_rd_0_Q_[63]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[7]\\\               : out   std_logic;
          \Z\\Fifo_rd_0_Q_[56]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[25]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[24]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[48]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[65]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[64]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[51]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[38]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[71]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[50]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[70]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[18]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[6]\\\               : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[71]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[70]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[69]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[68]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[67]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[66]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[65]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[64]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[63]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[62]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[61]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[60]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[59]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[58]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[57]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[56]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[55]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[54]\\\ : in    std_logic;
          \Z\\Fifo_rd_0_Q_[46]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[52]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[36]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[59]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[0]\\\               : out   std_logic;
          \Z\\Fifo_rd_0_Q_[16]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[57]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[41]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[53]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[40]\\\              : out   std_logic;
          Main_ctl4SD_0_fifo_rd                : in    std_logic;
          \Z\\Fifo_rd_0_Q_[31]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[28]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[30]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[42]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[11]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[10]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[55]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[68]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[54]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[49]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[9]\\\               : out   std_logic;
          \Z\\Fifo_rd_0_Q_[5]\\\               : out   std_logic;
          Fifo_rd_0_AFULL                      : out   std_logic;
          \Z\\Fifo_rd_0_Q_[32]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[47]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[43]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[12]\\\              : out   std_logic;
          Sdram_cmd_0_RFifo_we                 : in    std_logic;
          \Z\\Fifo_rd_0_Q_[26]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[39]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[19]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[37]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[3]\\\               : out   std_logic;
          \Z\\Fifo_rd_0_Q_[33]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[66]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[17]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[13]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[45]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[44]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[21]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[2]\\\               : out   std_logic;
          \Z\\Fifo_rd_0_Q_[20]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[61]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[35]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[34]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[60]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[15]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[14]\\\              : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[35]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[34]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[33]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[32]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[31]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[30]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[29]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[28]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[27]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[26]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[25]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[24]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[23]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[22]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[21]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[20]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[19]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[18]\\\ : in    std_logic;
          Main_ctl4SD_0_fifo_rst_n_0           : in    std_logic;
          \Z\\Fifo_rd_0_Q_[22]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[8]\\\               : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[53]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[52]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[51]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[50]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[49]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[48]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[47]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[46]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[45]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[44]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[43]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[42]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[41]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[40]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[39]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[38]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[37]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[36]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[17]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[16]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[15]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[14]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[13]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[12]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[11]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[10]\\\ : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[9]\\\  : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[8]\\\  : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[7]\\\  : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[6]\\\  : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[5]\\\  : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[4]\\\  : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[3]\\\  : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[2]\\\  : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[1]\\\  : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[0]\\\  : in    std_logic;
          Fifo_rd_1_VCC                        : in    std_logic;
          Main_ctl4SD_0_fifo_rst_n_3           : in    std_logic;
          \Z\\Fifo_rd_0_Q_[62]\\\              : out   std_logic;
          Main_ctl4SD_0_fifo_rst_n_1           : in    std_logic;
          \Z\\Fifo_rd_0_Q_[29]\\\              : out   std_logic;
          Main_ctl4SD_0_fifo_rst_n_2           : in    std_logic;
          PLL_Test1_0_Sys_66M_Clk              : in    std_logic;
          \Z\\Fifo_rd_0_Q_[58]\\\              : out   std_logic;
          Fifo_rd_1_GND                        : in    std_logic
        );

end Fifo_rd_1;

architecture DEF_ARCH of Fifo_rd_1 is 

  component INV
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XNOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component RAM512X18
    generic (MEMORYFILE:string := "");

    port( RADDR8 : in    std_logic := 'U';
          RADDR7 : in    std_logic := 'U';
          RADDR6 : in    std_logic := 'U';
          RADDR5 : in    std_logic := 'U';
          RADDR4 : in    std_logic := 'U';
          RADDR3 : in    std_logic := 'U';
          RADDR2 : in    std_logic := 'U';
          RADDR1 : in    std_logic := 'U';
          RADDR0 : in    std_logic := 'U';
          WADDR8 : in    std_logic := 'U';
          WADDR7 : in    std_logic := 'U';
          WADDR6 : in    std_logic := 'U';
          WADDR5 : in    std_logic := 'U';
          WADDR4 : in    std_logic := 'U';
          WADDR3 : in    std_logic := 'U';
          WADDR2 : in    std_logic := 'U';
          WADDR1 : in    std_logic := 'U';
          WADDR0 : in    std_logic := 'U';
          WD17   : in    std_logic := 'U';
          WD16   : in    std_logic := 'U';
          WD15   : in    std_logic := 'U';
          WD14   : in    std_logic := 'U';
          WD13   : in    std_logic := 'U';
          WD12   : in    std_logic := 'U';
          WD11   : in    std_logic := 'U';
          WD10   : in    std_logic := 'U';
          WD9    : in    std_logic := 'U';
          WD8    : in    std_logic := 'U';
          WD7    : in    std_logic := 'U';
          WD6    : in    std_logic := 'U';
          WD5    : in    std_logic := 'U';
          WD4    : in    std_logic := 'U';
          WD3    : in    std_logic := 'U';
          WD2    : in    std_logic := 'U';
          WD1    : in    std_logic := 'U';
          WD0    : in    std_logic := 'U';
          RW0    : in    std_logic := 'U';
          RW1    : in    std_logic := 'U';
          WW0    : in    std_logic := 'U';
          WW1    : in    std_logic := 'U';
          PIPE   : in    std_logic := 'U';
          REN    : in    std_logic := 'U';
          WEN    : in    std_logic := 'U';
          RCLK   : in    std_logic := 'U';
          WCLK   : in    std_logic := 'U';
          RESET  : in    std_logic := 'U';
          RD17   : out   std_logic;
          RD16   : out   std_logic;
          RD15   : out   std_logic;
          RD14   : out   std_logic;
          RD13   : out   std_logic;
          RD12   : out   std_logic;
          RD11   : out   std_logic;
          RD10   : out   std_logic;
          RD9    : out   std_logic;
          RD8    : out   std_logic;
          RD7    : out   std_logic;
          RD6    : out   std_logic;
          RD5    : out   std_logic;
          RD4    : out   std_logic;
          RD3    : out   std_logic;
          RD2    : out   std_logic;
          RD1    : out   std_logic;
          RD0    : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AND3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component NAND3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AO1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component BUFF
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NAND2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal DVLDI_2, DVLDI, DVLDI_1, DVLDI_0, AND2_25_Y, AND3_1_Y, 
        XNOR2_6_Y, AND2_28_Y, MEM_RADDR_0_net, MEMORYRE, 
        XNOR2_8_Y, MEM_RADDR_3_net, WBINNXTSHIFT_3_net, XOR2_36_Y, 
        MEM_RADDR_4_net, QXI_58_net, QXI_29_net, 
        RBINNXTSHIFT_2_net, XOR2_10_Y, AO1_8_Y, QXI_62_net, 
        QXI_0_net, QXI_1_net, QXI_2_net, QXI_3_net, QXI_4_net, 
        QXI_5_net, QXI_6_net, QXI_7_net, QXI_8_net, QXI_9_net, 
        QXI_10_net, QXI_11_net, QXI_12_net, QXI_13_net, 
        QXI_14_net, QXI_15_net, QXI_16_net, QXI_17_net, 
        MEM_RADDR_1_net, MEM_RADDR_2_net, MEMRENEG, 
        MEM_WADDR_0_net, MEM_WADDR_1_net, MEM_WADDR_2_net, 
        MEM_WADDR_3_net, MEMWENEG, AO1_4_Y, XOR2_11_Y, AO1_0_Y, 
        AND2_3_Y, NAND2_1_Y, DFN1P0_EMPTY_0, XOR2_0_Y, 
        WBINNXTSHIFT_1_net, AND2_8_Y, AND2_21_Y, QXI_36_net, 
        QXI_37_net, QXI_38_net, QXI_39_net, QXI_40_net, 
        QXI_41_net, QXI_42_net, QXI_43_net, QXI_44_net, 
        QXI_45_net, QXI_46_net, QXI_47_net, QXI_48_net, 
        QXI_49_net, QXI_50_net, QXI_51_net, QXI_52_net, 
        QXI_53_net, QXI_22_net, RBINNXTSHIFT_0_net, QXI_18_net, 
        QXI_19_net, QXI_20_net, QXI_21_net, QXI_23_net, 
        QXI_24_net, QXI_25_net, QXI_26_net, QXI_27_net, 
        QXI_28_net, QXI_30_net, QXI_31_net, QXI_32_net, 
        QXI_33_net, QXI_34_net, QXI_35_net, XOR2_28_Y, QXI_60_net, 
        RBINNXTSHIFT_1_net, XOR2_29_Y, QXI_61_net, XOR2_3_Y, 
        INV_2_Y, MEMORYWE, WDIFF_4_net, XOR2_21_Y, AO1_6_Y, 
        AO1_5_Y, AND2_24_Y, AO1_11_Y, XNOR2_5_Y, FULLINT, 
        AND2_7_Y, XOR2_23_Y, AND2_4_Y, XNOR2_7_Y, OR2A_0_Y, 
        WDIFF_2_net, AO1_13_Y, XOR2_4_Y, NOR2A_0_Y, 
        WBINNXTSHIFT_0_net, AND2_17_Y, INV_3_Y, QXI_66_net, 
        EMPTYINT, XOR2_35_Y, AO1_10_Y, AND2_1_Y, AOI1_0_Y, 
        AND2_6_Y, NAND3A_1_Y, NOR3_0_Y, OA1A_0_Y, WDIFF_3_net, 
        WDIFF_1_net, XOR2_14_Y, AND2A_0_Y, XOR2_2_Y, XOR2_18_Y, 
        AND2_18_Y, NAND2_0_Y, XNOR2_10_Y, RBINNXTSHIFT_4_net, 
        MEM_WADDR_4_net, AND2A_1_Y, DFN1C0_FULL_0, NOR3A_0_Y, 
        NAND3A_0_Y, OR2_0_Y, OR2A_1_Y, AO1C_0_Y, WDIFF_0_net, 
        AND2_9_Y, QXI_54_net, OR3_0_Y, AND2_22_Y, AND2_2_Y, 
        QXI_68_net, QXI_55_net, XOR2_32_Y, RBINNXTSHIFT_3_net, 
        AO1_7_Y, XNOR2_3_Y, INV_1_Y, XOR2_7_Y, WBINNXTSHIFT_2_net, 
        INV_4_Y, XNOR2_1_Y, AND2_13_Y, XOR2_9_Y, AO1_3_Y, 
        AND2_12_Y, QXI_57_net, XOR2_13_Y, QXI_59_net, XNOR2_4_Y, 
        XOR2_20_Y, OA1C_0_Y, WBINNXTSHIFT_4_net, XOR2_16_Y, 
        QXI_56_net, QXI_63_net, QXI_64_net, QXI_65_net, 
        QXI_67_net, QXI_69_net, QXI_70_net, QXI_71_net, AND2_31_Y, 
        XNOR2_0_Y, XOR2_1_Y, XNOR2_2_Y, AND3_0_Y, XNOR2_9_Y, 
        INV_0_Y, \GND\, \VCC\, GND_0, VCC_0 : std_logic;

begin 


    INV_0 : INV
      port map(A => MEM_RADDR_4_net, Y => INV_0_Y);
    
    NOR3_0 : NOR3
      port map(A => OA1A_0_Y, B => AND2A_0_Y, C => OA1C_0_Y, Y
         => NOR3_0_Y);
    
    AND2_2 : AND2
      port map(A => INV_1_Y, B => INV_3_Y, Y => AND2_2_Y);
    
    DFN1E1C0_Q_27_inst : DFN1E1C0
      port map(D => QXI_27_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_1, E => DVLDI_0, Q => 
        \Z\\Fifo_rd_0_Q_[27]\\\);
    
    AO1_11 : AO1
      port map(A => XOR2_1_Y, B => AND2_4_Y, C => AND2_21_Y, Y
         => AO1_11_Y);
    
    AND2_22 : AND2
      port map(A => WBINNXTSHIFT_1_net, B => INV_1_Y, Y => 
        AND2_22_Y);
    
    XNOR2_9 : XNOR2
      port map(A => MEM_RADDR_2_net, B => WBINNXTSHIFT_2_net, Y
         => XNOR2_9_Y);
    
    DFN1C0_FULL : DFN1C0
      port map(D => FULLINT, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => Main_ctl4SD_0_fifo_rst_n_0, Q => DFN1C0_FULL_0);
    
    DFN1E1C0_Q_37_inst : DFN1E1C0
      port map(D => QXI_37_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_1, E => DVLDI_1, Q => 
        \Z\\Fifo_rd_0_Q_[37]\\\);
    
    DFN1E1C0_Q_23_inst : DFN1E1C0
      port map(D => QXI_23_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_1, E => DVLDI_0, Q => 
        \Z\\Fifo_rd_0_Q_[23]\\\);
    
    XOR2_23 : XOR2
      port map(A => MEM_RADDR_4_net, B => WBINNXTSHIFT_4_net, Y
         => XOR2_23_Y);
    
    XOR2_1 : XOR2
      port map(A => MEM_RADDR_3_net, B => Fifo_rd_1_GND, Y => 
        XOR2_1_Y);
    
    DFN1E1C0_Q_54_inst : DFN1E1C0
      port map(D => QXI_54_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_2, E => DVLDI_2, Q => 
        \Z\\Fifo_rd_0_Q_[54]\\\);
    
    DFN1E1C0_Q_33_inst : DFN1E1C0
      port map(D => QXI_33_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_1, E => DVLDI_1, Q => 
        \Z\\Fifo_rd_0_Q_[33]\\\);
    
    INV_1 : INV
      port map(A => MEM_RADDR_1_net, Y => INV_1_Y);
    
    AO1_7 : AO1
      port map(A => XOR2_7_Y, B => OR3_0_Y, C => AND2_31_Y, Y => 
        AO1_7_Y);
    
    AND2_18 : AND2
      port map(A => MEM_WADDR_1_net, B => Fifo_rd_1_GND, Y => 
        AND2_18_Y);
    
    DFN1C0_MEM_WADDR_2_inst : DFN1C0
      port map(D => WBINNXTSHIFT_2_net, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => 
        Main_ctl4SD_0_fifo_rst_n_0, Q => MEM_WADDR_2_net);
    
    AND2_1 : AND2
      port map(A => MEM_WADDR_3_net, B => Fifo_rd_1_GND, Y => 
        AND2_1_Y);
    
    AO1_8 : AO1
      port map(A => XOR2_2_Y, B => AND2_28_Y, C => AND2_13_Y, Y
         => AO1_8_Y);
    
    DFN1E1C0_Q_61_inst : DFN1E1C0
      port map(D => QXI_61_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_3, E => DVLDI_2, Q => 
        \Z\\Fifo_rd_0_Q_[61]\\\);
    
    XOR2_20 : XOR2
      port map(A => WBINNXTSHIFT_2_net, B => INV_4_Y, Y => 
        XOR2_20_Y);
    
    DFN1E1C0_Q_2_inst : DFN1E1C0
      port map(D => QXI_2_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_1, E => DVLDI_0, Q => 
        \Z\\Fifo_rd_0_Q_[2]\\\);
    
    AND2_7 : AND2
      port map(A => AND3_0_Y, B => XNOR2_8_Y, Y => AND2_7_Y);
    
    AND2_12 : AND2
      port map(A => XOR2_11_Y, B => XOR2_35_Y, Y => AND2_12_Y);
    
    AND2A_1 : AND2A
      port map(A => DFN1P0_EMPTY_0, B => Main_ctl4SD_0_fifo_rd, Y
         => AND2A_1_Y);
    
    DFN1E1C0_Q_65_inst : DFN1E1C0
      port map(D => QXI_65_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_3, E => DVLDI_2, Q => 
        \Z\\Fifo_rd_0_Q_[65]\\\);
    
    AND2_EMPTYINT : AND2
      port map(A => AND2_25_Y, B => XNOR2_10_Y, Y => EMPTYINT);
    
    RAM512X18_QXI_17_inst : RAM512X18
      port map(RADDR8 => Fifo_rd_1_GND, RADDR7 => Fifo_rd_1_GND, 
        RADDR6 => Fifo_rd_1_GND, RADDR5 => Fifo_rd_1_GND, RADDR4
         => Fifo_rd_1_GND, RADDR3 => MEM_RADDR_3_net, RADDR2 => 
        MEM_RADDR_2_net, RADDR1 => MEM_RADDR_1_net, RADDR0 => 
        MEM_RADDR_0_net, WADDR8 => Fifo_rd_1_GND, WADDR7 => 
        Fifo_rd_1_GND, WADDR6 => Fifo_rd_1_GND, WADDR5 => 
        Fifo_rd_1_GND, WADDR4 => Fifo_rd_1_GND, WADDR3 => 
        MEM_WADDR_3_net, WADDR2 => MEM_WADDR_2_net, WADDR1 => 
        MEM_WADDR_1_net, WADDR0 => MEM_WADDR_0_net, WD17 => 
        \Z\\Sdram_data_0_Sys_dataOut_[17]\\\, WD16 => 
        \Z\\Sdram_data_0_Sys_dataOut_[16]\\\, WD15 => 
        \Z\\Sdram_data_0_Sys_dataOut_[15]\\\, WD14 => 
        \Z\\Sdram_data_0_Sys_dataOut_[14]\\\, WD13 => 
        \Z\\Sdram_data_0_Sys_dataOut_[13]\\\, WD12 => 
        \Z\\Sdram_data_0_Sys_dataOut_[12]\\\, WD11 => 
        \Z\\Sdram_data_0_Sys_dataOut_[11]\\\, WD10 => 
        \Z\\Sdram_data_0_Sys_dataOut_[10]\\\, WD9 => 
        \Z\\Sdram_data_0_Sys_dataOut_[9]\\\, WD8 => 
        \Z\\Sdram_data_0_Sys_dataOut_[8]\\\, WD7 => 
        \Z\\Sdram_data_0_Sys_dataOut_[7]\\\, WD6 => 
        \Z\\Sdram_data_0_Sys_dataOut_[6]\\\, WD5 => 
        \Z\\Sdram_data_0_Sys_dataOut_[5]\\\, WD4 => 
        \Z\\Sdram_data_0_Sys_dataOut_[4]\\\, WD3 => 
        \Z\\Sdram_data_0_Sys_dataOut_[3]\\\, WD2 => 
        \Z\\Sdram_data_0_Sys_dataOut_[2]\\\, WD1 => 
        \Z\\Sdram_data_0_Sys_dataOut_[1]\\\, WD0 => 
        \Z\\Sdram_data_0_Sys_dataOut_[0]\\\, RW0 => Fifo_rd_1_GND, 
        RW1 => Fifo_rd_1_VCC, WW0 => Fifo_rd_1_GND, WW1 => 
        Fifo_rd_1_VCC, PIPE => Fifo_rd_1_GND, REN => MEMRENEG, 
        WEN => MEMWENEG, RCLK => PLL_Test1_0_Sys_66M_Clk, WCLK
         => PLL_Test1_0_Sys_66M_Clk, RESET => 
        Main_ctl4SD_0_fifo_rst_n_3, RD17 => QXI_17_net, RD16 => 
        QXI_16_net, RD15 => QXI_15_net, RD14 => QXI_14_net, RD13
         => QXI_13_net, RD12 => QXI_12_net, RD11 => QXI_11_net, 
        RD10 => QXI_10_net, RD9 => QXI_9_net, RD8 => QXI_8_net, 
        RD7 => QXI_7_net, RD6 => QXI_6_net, RD5 => QXI_5_net, RD4
         => QXI_4_net, RD3 => QXI_3_net, RD2 => QXI_2_net, RD1
         => QXI_1_net, RD0 => QXI_0_net);
    
    XOR2_21 : XOR2
      port map(A => WBINNXTSHIFT_4_net, B => INV_0_Y, Y => 
        XOR2_21_Y);
    
    DFN1C0_MEM_RADDR_0_inst : DFN1C0
      port map(D => RBINNXTSHIFT_0_net, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => 
        Main_ctl4SD_0_fifo_rst_n_0, Q => MEM_RADDR_0_net);
    
    DFN1E1C0_Q_5_inst : DFN1E1C0
      port map(D => QXI_5_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_2, E => DVLDI_2, Q => 
        \Z\\Fifo_rd_0_Q_[5]\\\);
    
    DFN1E1C0_Q_14_inst : DFN1E1C0
      port map(D => QXI_14_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_0, E => DVLDI_0, Q => 
        \Z\\Fifo_rd_0_Q_[14]\\\);
    
    XOR2_16 : XOR2
      port map(A => MEM_WADDR_4_net, B => Fifo_rd_1_GND, Y => 
        XOR2_16_Y);
    
    DFN1E1C0_Q_66_inst : DFN1E1C0
      port map(D => QXI_66_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_3, E => DVLDI_2, Q => 
        \Z\\Fifo_rd_0_Q_[66]\\\);
    
    RAM512X18_QXI_53_inst : RAM512X18
      port map(RADDR8 => Fifo_rd_1_GND, RADDR7 => Fifo_rd_1_GND, 
        RADDR6 => Fifo_rd_1_GND, RADDR5 => Fifo_rd_1_GND, RADDR4
         => Fifo_rd_1_GND, RADDR3 => MEM_RADDR_3_net, RADDR2 => 
        MEM_RADDR_2_net, RADDR1 => MEM_RADDR_1_net, RADDR0 => 
        MEM_RADDR_0_net, WADDR8 => Fifo_rd_1_GND, WADDR7 => 
        Fifo_rd_1_GND, WADDR6 => Fifo_rd_1_GND, WADDR5 => 
        Fifo_rd_1_GND, WADDR4 => Fifo_rd_1_GND, WADDR3 => 
        MEM_WADDR_3_net, WADDR2 => MEM_WADDR_2_net, WADDR1 => 
        MEM_WADDR_1_net, WADDR0 => MEM_WADDR_0_net, WD17 => 
        \Z\\Sdram_data_0_Sys_dataOut_[53]\\\, WD16 => 
        \Z\\Sdram_data_0_Sys_dataOut_[52]\\\, WD15 => 
        \Z\\Sdram_data_0_Sys_dataOut_[51]\\\, WD14 => 
        \Z\\Sdram_data_0_Sys_dataOut_[50]\\\, WD13 => 
        \Z\\Sdram_data_0_Sys_dataOut_[49]\\\, WD12 => 
        \Z\\Sdram_data_0_Sys_dataOut_[48]\\\, WD11 => 
        \Z\\Sdram_data_0_Sys_dataOut_[47]\\\, WD10 => 
        \Z\\Sdram_data_0_Sys_dataOut_[46]\\\, WD9 => 
        \Z\\Sdram_data_0_Sys_dataOut_[45]\\\, WD8 => 
        \Z\\Sdram_data_0_Sys_dataOut_[44]\\\, WD7 => 
        \Z\\Sdram_data_0_Sys_dataOut_[43]\\\, WD6 => 
        \Z\\Sdram_data_0_Sys_dataOut_[42]\\\, WD5 => 
        \Z\\Sdram_data_0_Sys_dataOut_[41]\\\, WD4 => 
        \Z\\Sdram_data_0_Sys_dataOut_[40]\\\, WD3 => 
        \Z\\Sdram_data_0_Sys_dataOut_[39]\\\, WD2 => 
        \Z\\Sdram_data_0_Sys_dataOut_[38]\\\, WD1 => 
        \Z\\Sdram_data_0_Sys_dataOut_[37]\\\, WD0 => 
        \Z\\Sdram_data_0_Sys_dataOut_[36]\\\, RW0 => 
        Fifo_rd_1_GND, RW1 => Fifo_rd_1_VCC, WW0 => Fifo_rd_1_GND, 
        WW1 => Fifo_rd_1_VCC, PIPE => Fifo_rd_1_GND, REN => 
        MEMRENEG, WEN => MEMWENEG, RCLK => 
        PLL_Test1_0_Sys_66M_Clk, WCLK => PLL_Test1_0_Sys_66M_Clk, 
        RESET => Main_ctl4SD_0_fifo_rst_n_3, RD17 => QXI_53_net, 
        RD16 => QXI_52_net, RD15 => QXI_51_net, RD14 => 
        QXI_50_net, RD13 => QXI_49_net, RD12 => QXI_48_net, RD11
         => QXI_47_net, RD10 => QXI_46_net, RD9 => QXI_45_net, 
        RD8 => QXI_44_net, RD7 => QXI_43_net, RD6 => QXI_42_net, 
        RD5 => QXI_41_net, RD4 => QXI_40_net, RD3 => QXI_39_net, 
        RD2 => QXI_38_net, RD1 => QXI_37_net, RD0 => QXI_36_net);
    
    DFN1E1C0_Q_62_inst : DFN1E1C0
      port map(D => QXI_62_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_3, E => DVLDI_2, Q => 
        \Z\\Fifo_rd_0_Q_[62]\\\);
    
    OR2_0 : OR2
      port map(A => AOI1_0_Y, B => DFN1C0_FULL_0, Y => OR2_0_Y);
    
    MEMWEBUBBLE : INV
      port map(A => MEMORYWE, Y => MEMWENEG);
    
    AND2_6 : AND2
      port map(A => XNOR2_4_Y, B => XNOR2_1_Y, Y => AND2_6_Y);
    
    AND3_0 : AND3
      port map(A => XNOR2_0_Y, B => XNOR2_7_Y, C => XNOR2_9_Y, Y
         => AND3_0_Y);
    
    DFN1E1C0_Q_0_inst : DFN1E1C0
      port map(D => QXI_0_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_0, E => DVLDI_0, Q => 
        \Z\\Fifo_rd_0_Q_[0]\\\);
    
    INV_3 : INV
      port map(A => NOR2A_0_Y, Y => INV_3_Y);
    
    XNOR2_2 : XNOR2
      port map(A => RBINNXTSHIFT_1_net, B => MEM_WADDR_1_net, Y
         => XNOR2_2_Y);
    
    DFN1E1C0_Q_29_inst : DFN1E1C0
      port map(D => QXI_29_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_1, E => DVLDI_0, Q => 
        \Z\\Fifo_rd_0_Q_[29]\\\);
    
    XOR2_WBINNXTSHIFT_2_inst : XOR2
      port map(A => XOR2_13_Y, B => AO1_0_Y, Y => 
        WBINNXTSHIFT_2_net);
    
    XOR2_4 : XOR2
      port map(A => MEM_RADDR_2_net, B => Fifo_rd_1_GND, Y => 
        XOR2_4_Y);
    
    AND3_1 : AND3
      port map(A => XNOR2_3_Y, B => XNOR2_2_Y, C => XNOR2_5_Y, Y
         => AND3_1_Y);
    
    AND2_24 : AND2
      port map(A => XOR2_4_Y, B => XOR2_1_Y, Y => AND2_24_Y);
    
    XNOR2_0 : XNOR2
      port map(A => MEM_RADDR_0_net, B => WBINNXTSHIFT_0_net, Y
         => XNOR2_0_Y);
    
    DFN1E1C0_Q_39_inst : DFN1E1C0
      port map(D => QXI_39_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_1, E => DVLDI_1, Q => 
        \Z\\Fifo_rd_0_Q_[39]\\\);
    
    AND2_31 : AND2
      port map(A => WBINNXTSHIFT_2_net, B => INV_4_Y, Y => 
        AND2_31_Y);
    
    GND_i : GND
      port map(Y => \GND\);
    
    XOR2_WBINNXTSHIFT_0_inst : XOR2
      port map(A => MEM_WADDR_0_net, B => MEMORYWE, Y => 
        WBINNXTSHIFT_0_net);
    
    XOR2_18 : XOR2
      port map(A => MEM_WADDR_1_net, B => Fifo_rd_1_GND, Y => 
        XOR2_18_Y);
    
    DFN1E1C0_Q_41_inst : DFN1E1C0
      port map(D => QXI_41_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_2, E => DVLDI_1, Q => 
        \Z\\Fifo_rd_0_Q_[41]\\\);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    NAND3A_0 : NAND3A
      port map(A => WDIFF_1_net, B => Fifo_rd_1_GND, C => 
        OR2A_1_Y, Y => NAND3A_0_Y);
    
    DFN1E1C0_Q_45_inst : DFN1E1C0
      port map(D => QXI_45_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_2, E => DVLDI_1, Q => 
        \Z\\Fifo_rd_0_Q_[45]\\\);
    
    XOR2_RBINNXTSHIFT_2_inst : XOR2
      port map(A => XOR2_10_Y, B => AO1_8_Y, Y => 
        RBINNXTSHIFT_2_net);
    
    DFN1E1C0_Q_67_inst : DFN1E1C0
      port map(D => QXI_67_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_3, E => DVLDI_2, Q => 
        \Z\\Fifo_rd_0_Q_[67]\\\);
    
    MEMREBUBBLE : INV
      port map(A => MEMORYRE, Y => MEMRENEG);
    
    DFN1E1C0_Q_20_inst : DFN1E1C0
      port map(D => QXI_20_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_1, E => DVLDI_0, Q => 
        \Z\\Fifo_rd_0_Q_[20]\\\);
    
    DFN1E1C0_Q_63_inst : DFN1E1C0
      port map(D => QXI_63_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_3, E => DVLDI_2, Q => 
        \Z\\Fifo_rd_0_Q_[63]\\\);
    
    XOR2_RBINNXTSHIFT_0_inst : XOR2
      port map(A => MEM_RADDR_0_net, B => MEMORYRE, Y => 
        RBINNXTSHIFT_0_net);
    
    XOR2_WBINNXTSHIFT_1_inst : XOR2
      port map(A => XOR2_0_Y, B => AND2_8_Y, Y => 
        WBINNXTSHIFT_1_net);
    
    DFN1E1C0_Q_30_inst : DFN1E1C0
      port map(D => QXI_30_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_1, E => DVLDI_0, Q => 
        \Z\\Fifo_rd_0_Q_[30]\\\);
    
    AND2_3 : AND2
      port map(A => MEM_WADDR_2_net, B => Fifo_rd_1_GND, Y => 
        AND2_3_Y);
    
    DFN1E1C0_Q_28_inst : DFN1E1C0
      port map(D => QXI_28_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_1, E => DVLDI_0, Q => 
        \Z\\Fifo_rd_0_Q_[28]\\\);
    
    DFN1E1C0_Q_46_inst : DFN1E1C0
      port map(D => QXI_46_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_2, E => DVLDI_1, Q => 
        \Z\\Fifo_rd_0_Q_[46]\\\);
    
    XNOR2_6 : XNOR2
      port map(A => RBINNXTSHIFT_3_net, B => MEM_WADDR_3_net, Y
         => XNOR2_6_Y);
    
    OA1C_0 : OA1C
      port map(A => Fifo_rd_1_VCC, B => WDIFF_3_net, C => 
        Fifo_rd_1_GND, Y => OA1C_0_Y);
    
    INV_4 : INV
      port map(A => MEM_RADDR_2_net, Y => INV_4_Y);
    
    OR2A_1 : OR2A
      port map(A => WDIFF_2_net, B => Fifo_rd_1_GND, Y => 
        OR2A_1_Y);
    
    DFN1E1C0_Q_38_inst : DFN1E1C0
      port map(D => QXI_38_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_1, E => DVLDI_1, Q => 
        \Z\\Fifo_rd_0_Q_[38]\\\);
    
    DFN1E1C0_Q_42_inst : DFN1E1C0
      port map(D => QXI_42_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_2, E => DVLDI_1, Q => 
        \Z\\Fifo_rd_0_Q_[42]\\\);
    
    DFN1E1C0_Q_51_inst : DFN1E1C0
      port map(D => QXI_51_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_2, E => DVLDI_1, Q => 
        \Z\\Fifo_rd_0_Q_[51]\\\);
    
    XOR2_9 : XOR2
      port map(A => WBINNXTSHIFT_3_net, B => INV_2_Y, Y => 
        XOR2_9_Y);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    XOR2_RBINNXTSHIFT_1_inst : XOR2
      port map(A => XOR2_29_Y, B => AND2_28_Y, Y => 
        RBINNXTSHIFT_1_net);
    
    XNOR2_4 : XNOR2
      port map(A => Fifo_rd_1_VCC, B => WDIFF_3_net, Y => 
        XNOR2_4_Y);
    
    DFN1E1C0_Q_55_inst : DFN1E1C0
      port map(D => QXI_55_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_2, E => DVLDI_2, Q => 
        \Z\\Fifo_rd_0_Q_[55]\\\);
    
    DFN1E1C0_Q_1_inst : DFN1E1C0
      port map(D => QXI_1_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_1, E => DVLDI_0, Q => 
        \Z\\Fifo_rd_0_Q_[1]\\\);
    
    DFN1C0_MEM_WADDR_4_inst : DFN1C0
      port map(D => WBINNXTSHIFT_4_net, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => 
        Main_ctl4SD_0_fifo_rst_n_0, Q => MEM_WADDR_4_net);
    
    DFN1E1C0_Q_4_inst : DFN1E1C0
      port map(D => QXI_4_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_2, E => DVLDI_1, Q => 
        \Z\\Fifo_rd_0_Q_[4]\\\);
    
    XOR2_13 : XOR2
      port map(A => MEM_WADDR_2_net, B => Fifo_rd_1_GND, Y => 
        XOR2_13_Y);
    
    DFN1E1C0_Q_8_inst : DFN1E1C0
      port map(D => QXI_8_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_3, E => DVLDI_2, Q => 
        \Z\\Fifo_rd_0_Q_[8]\\\);
    
    XOR2_WBINNXTSHIFT_3_inst : XOR2
      port map(A => XOR2_32_Y, B => AO1_4_Y, Y => 
        WBINNXTSHIFT_3_net);
    
    XOR2_WDIFF_4_inst : XOR2
      port map(A => XOR2_21_Y, B => AO1_6_Y, Y => WDIFF_4_net);
    
    DFN1E1C0_Q_56_inst : DFN1E1C0
      port map(D => QXI_56_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_2, E => DVLDI_2, Q => 
        \Z\\Fifo_rd_0_Q_[56]\\\);
    
    AO1_3 : AO1
      port map(A => AND2_12_Y, B => AO1_0_Y, C => AO1_10_Y, Y => 
        AO1_3_Y);
    
    DFN1E1C0_Q_70_inst : DFN1E1C0
      port map(D => QXI_70_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_3, E => DVLDI_2, Q => 
        \Z\\Fifo_rd_0_Q_[70]\\\);
    
    DFN1E1C0_Q_47_inst : DFN1E1C0
      port map(D => QXI_47_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_2, E => DVLDI_1, Q => 
        \Z\\Fifo_rd_0_Q_[47]\\\);
    
    DFN1E1C0_Q_52_inst : DFN1E1C0
      port map(D => QXI_52_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_2, E => DVLDI_1, Q => 
        \Z\\Fifo_rd_0_Q_[52]\\\);
    
    AO1C_0 : AO1C
      port map(A => Fifo_rd_1_GND, B => WDIFF_1_net, C => 
        Fifo_rd_1_GND, Y => AO1C_0_Y);
    
    DFN1E1C0_Q_7_inst : DFN1E1C0
      port map(D => QXI_7_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_3, E => DVLDI_2, Q => 
        \Z\\Fifo_rd_0_Q_[7]\\\);
    
    DFN1E1C0_Q_43_inst : DFN1E1C0
      port map(D => QXI_43_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_2, E => DVLDI_1, Q => 
        \Z\\Fifo_rd_0_Q_[43]\\\);
    
    AND2_13 : AND2
      port map(A => MEM_RADDR_1_net, B => Fifo_rd_1_GND, Y => 
        AND2_13_Y);
    
    DFN1E1C0_Q_11_inst : DFN1E1C0
      port map(D => QXI_11_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_0, E => DVLDI_0, Q => 
        \Z\\Fifo_rd_0_Q_[11]\\\);
    
    DFN1C0_DVLDI_RNI2T66 : BUFF
      port map(A => DVLDI, Y => DVLDI_1);
    
    XOR2_10 : XOR2
      port map(A => MEM_RADDR_2_net, B => Fifo_rd_1_GND, Y => 
        XOR2_10_Y);
    
    XNOR2_1 : XNOR2
      port map(A => Fifo_rd_1_GND, B => WDIFF_4_net, Y => 
        XNOR2_1_Y);
    
    XOR2_RBINNXTSHIFT_3_inst : XOR2
      port map(A => XOR2_28_Y, B => AO1_13_Y, Y => 
        RBINNXTSHIFT_3_net);
    
    DFN1E1C0_Q_15_inst : DFN1E1C0
      port map(D => QXI_15_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_0, E => DVLDI_0, Q => 
        \Z\\Fifo_rd_0_Q_[15]\\\);
    
    DFN1E1C0_Q_69_inst : DFN1E1C0
      port map(D => QXI_69_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_3, E => DVLDI_2, Q => 
        \Z\\Fifo_rd_0_Q_[69]\\\);
    
    AND2_MEMORYRE : AND2
      port map(A => NAND2_1_Y, B => Main_ctl4SD_0_fifo_rd, Y => 
        MEMORYRE);
    
    XOR2_7 : XOR2
      port map(A => WBINNXTSHIFT_2_net, B => INV_4_Y, Y => 
        XOR2_7_Y);
    
    XOR2_14 : XOR2
      port map(A => WBINNXTSHIFT_1_net, B => INV_1_Y, Y => 
        XOR2_14_Y);
    
    XOR2_11 : XOR2
      port map(A => MEM_WADDR_2_net, B => Fifo_rd_1_GND, Y => 
        XOR2_11_Y);
    
    XNOR2_3 : XNOR2
      port map(A => RBINNXTSHIFT_0_net, B => MEM_WADDR_0_net, Y
         => XNOR2_3_Y);
    
    DFN1E1C0_Q_24_inst : DFN1E1C0
      port map(D => QXI_24_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_1, E => DVLDI_0, Q => 
        \Z\\Fifo_rd_0_Q_[24]\\\);
    
    DFN1E1C0_Q_34_inst : DFN1E1C0
      port map(D => QXI_34_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_1, E => DVLDI_1, Q => 
        \Z\\Fifo_rd_0_Q_[34]\\\);
    
    DFN1E1C0_Q_57_inst : DFN1E1C0
      port map(D => QXI_57_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_2, E => DVLDI_2, Q => 
        \Z\\Fifo_rd_0_Q_[57]\\\);
    
    DFN1E1C0_Q_16_inst : DFN1E1C0
      port map(D => QXI_16_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_0, E => DVLDI_0, Q => 
        \Z\\Fifo_rd_0_Q_[16]\\\);
    
    DFN1C0_MEM_RADDR_3_inst : DFN1C0
      port map(D => RBINNXTSHIFT_3_net, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => 
        Main_ctl4SD_0_fifo_rst_n_0, Q => MEM_RADDR_3_net);
    
    AO1_6 : AO1
      port map(A => XOR2_3_Y, B => AO1_7_Y, C => AND2_9_Y, Y => 
        AO1_6_Y);
    
    DFN1E1C0_Q_12_inst : DFN1E1C0
      port map(D => QXI_12_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_0, E => DVLDI_0, Q => 
        \Z\\Fifo_rd_0_Q_[12]\\\);
    
    DFN1E1C0_Q_53_inst : DFN1E1C0
      port map(D => QXI_53_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_2, E => DVLDI_2, Q => 
        \Z\\Fifo_rd_0_Q_[53]\\\);
    
    XOR2_WBINNXTSHIFT_4_inst : XOR2
      port map(A => XOR2_16_Y, B => AO1_3_Y, Y => 
        WBINNXTSHIFT_4_net);
    
    DFN1E1C0_Q_60_inst : DFN1E1C0
      port map(D => QXI_60_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_3, E => DVLDI_2, Q => 
        \Z\\Fifo_rd_0_Q_[60]\\\);
    
    XOR2_32 : XOR2
      port map(A => MEM_WADDR_3_net, B => Fifo_rd_1_GND, Y => 
        XOR2_32_Y);
    
    OR3_0 : OR3
      port map(A => AND2_22_Y, B => AND2_17_Y, C => AND2_2_Y, Y
         => OR3_0_Y);
    
    AND2_9 : AND2
      port map(A => WBINNXTSHIFT_3_net, B => INV_2_Y, Y => 
        AND2_9_Y);
    
    RAM512X18_QXI_71_inst : RAM512X18
      port map(RADDR8 => Fifo_rd_1_GND, RADDR7 => Fifo_rd_1_GND, 
        RADDR6 => Fifo_rd_1_GND, RADDR5 => Fifo_rd_1_GND, RADDR4
         => Fifo_rd_1_GND, RADDR3 => MEM_RADDR_3_net, RADDR2 => 
        MEM_RADDR_2_net, RADDR1 => MEM_RADDR_1_net, RADDR0 => 
        MEM_RADDR_0_net, WADDR8 => Fifo_rd_1_GND, WADDR7 => 
        Fifo_rd_1_GND, WADDR6 => Fifo_rd_1_GND, WADDR5 => 
        Fifo_rd_1_GND, WADDR4 => Fifo_rd_1_GND, WADDR3 => 
        MEM_WADDR_3_net, WADDR2 => MEM_WADDR_2_net, WADDR1 => 
        MEM_WADDR_1_net, WADDR0 => MEM_WADDR_0_net, WD17 => 
        \Z\\Sdram_data_0_Sys_dataOut_[71]\\\, WD16 => 
        \Z\\Sdram_data_0_Sys_dataOut_[70]\\\, WD15 => 
        \Z\\Sdram_data_0_Sys_dataOut_[69]\\\, WD14 => 
        \Z\\Sdram_data_0_Sys_dataOut_[68]\\\, WD13 => 
        \Z\\Sdram_data_0_Sys_dataOut_[67]\\\, WD12 => 
        \Z\\Sdram_data_0_Sys_dataOut_[66]\\\, WD11 => 
        \Z\\Sdram_data_0_Sys_dataOut_[65]\\\, WD10 => 
        \Z\\Sdram_data_0_Sys_dataOut_[64]\\\, WD9 => 
        \Z\\Sdram_data_0_Sys_dataOut_[63]\\\, WD8 => 
        \Z\\Sdram_data_0_Sys_dataOut_[62]\\\, WD7 => 
        \Z\\Sdram_data_0_Sys_dataOut_[61]\\\, WD6 => 
        \Z\\Sdram_data_0_Sys_dataOut_[60]\\\, WD5 => 
        \Z\\Sdram_data_0_Sys_dataOut_[59]\\\, WD4 => 
        \Z\\Sdram_data_0_Sys_dataOut_[58]\\\, WD3 => 
        \Z\\Sdram_data_0_Sys_dataOut_[57]\\\, WD2 => 
        \Z\\Sdram_data_0_Sys_dataOut_[56]\\\, WD1 => 
        \Z\\Sdram_data_0_Sys_dataOut_[55]\\\, WD0 => 
        \Z\\Sdram_data_0_Sys_dataOut_[54]\\\, RW0 => 
        Fifo_rd_1_GND, RW1 => Fifo_rd_1_VCC, WW0 => Fifo_rd_1_GND, 
        WW1 => Fifo_rd_1_VCC, PIPE => Fifo_rd_1_GND, REN => 
        MEMRENEG, WEN => MEMWENEG, RCLK => 
        PLL_Test1_0_Sys_66M_Clk, WCLK => PLL_Test1_0_Sys_66M_Clk, 
        RESET => Main_ctl4SD_0_fifo_rst_n_3, RD17 => QXI_71_net, 
        RD16 => QXI_70_net, RD15 => QXI_69_net, RD14 => 
        QXI_68_net, RD13 => QXI_67_net, RD12 => QXI_66_net, RD11
         => QXI_65_net, RD10 => QXI_64_net, RD9 => QXI_63_net, 
        RD8 => QXI_62_net, RD7 => QXI_61_net, RD6 => QXI_60_net, 
        RD5 => QXI_59_net, RD4 => QXI_58_net, RD3 => QXI_57_net, 
        RD2 => QXI_56_net, RD1 => QXI_55_net, RD0 => QXI_54_net);
    
    NOR3A_0 : NOR3A
      port map(A => OR2A_1_Y, B => AO1C_0_Y, C => WDIFF_0_net, Y
         => NOR3A_0_Y);
    
    DFN1E1C0_Q_68_inst : DFN1E1C0
      port map(D => QXI_68_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_3, E => DVLDI_2, Q => 
        \Z\\Fifo_rd_0_Q_[68]\\\);
    
    DFN1C0_AFULL : DFN1C0
      port map(D => OR2_0_Y, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => Main_ctl4SD_0_fifo_rst_n_0, Q => Fifo_rd_0_AFULL);
    
    INV_2 : INV
      port map(A => MEM_RADDR_3_net, Y => INV_2_Y);
    
    DFN1C0_MEM_WADDR_1_inst : DFN1C0
      port map(D => WBINNXTSHIFT_1_net, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => 
        Main_ctl4SD_0_fifo_rst_n_0, Q => MEM_WADDR_1_net);
    
    NAND3A_1 : NAND3A
      port map(A => NOR3A_0_Y, B => OR2A_0_Y, C => NAND3A_0_Y, Y
         => NAND3A_1_Y);
    
    NAND2_0 : NAND2
      port map(A => DFN1C0_FULL_0, B => Fifo_rd_1_VCC, Y => 
        NAND2_0_Y);
    
    DFN1E1C0_Q_3_inst : DFN1E1C0
      port map(D => QXI_3_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_2, E => DVLDI_1, Q => 
        \Z\\Fifo_rd_0_Q_[3]\\\);
    
    XOR2_RBINNXTSHIFT_4_inst : XOR2
      port map(A => XOR2_36_Y, B => AO1_5_Y, Y => 
        RBINNXTSHIFT_4_net);
    
    DFN1C0_DVLDI : DFN1C0
      port map(D => AND2A_1_Y, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_0, Q => DVLDI);
    
    XNOR2_10 : XNOR2
      port map(A => RBINNXTSHIFT_4_net, B => MEM_WADDR_4_net, Y
         => XNOR2_10_Y);
    
    AND2_MEMORYWE : AND2
      port map(A => NAND2_0_Y, B => Sdram_cmd_0_RFifo_we, Y => 
        MEMORYWE);
    
    DFN1E1C0_Q_49_inst : DFN1E1C0
      port map(D => QXI_49_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_2, E => DVLDI_1, Q => 
        \Z\\Fifo_rd_0_Q_[49]\\\);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    DFN1E1C0_Q_17_inst : DFN1E1C0
      port map(D => QXI_17_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_0, E => DVLDI_0, Q => 
        \Z\\Fifo_rd_0_Q_[17]\\\);
    
    AO1_0 : AO1
      port map(A => XOR2_18_Y, B => AND2_8_Y, C => AND2_18_Y, Y
         => AO1_0_Y);
    
    XOR2_29 : XOR2
      port map(A => MEM_RADDR_1_net, B => Fifo_rd_1_GND, Y => 
        XOR2_29_Y);
    
    DFN1C0_DVLDI_RNI2T66_1 : BUFF
      port map(A => DVLDI, Y => DVLDI_2);
    
    XOR2_2 : XOR2
      port map(A => MEM_RADDR_1_net, B => Fifo_rd_1_GND, Y => 
        XOR2_2_Y);
    
    DFN1C0_MEM_WADDR_0_inst : DFN1C0
      port map(D => WBINNXTSHIFT_0_net, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => 
        Main_ctl4SD_0_fifo_rst_n_0, Q => MEM_WADDR_0_net);
    
    DFN1E1C0_Q_13_inst : DFN1E1C0
      port map(D => QXI_13_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_0, E => DVLDI_0, Q => 
        \Z\\Fifo_rd_0_Q_[13]\\\);
    
    AND2A_0 : AND2A
      port map(A => Fifo_rd_1_GND, B => WDIFF_4_net, Y => 
        AND2A_0_Y);
    
    OA1A_0 : OA1A
      port map(A => Fifo_rd_1_VCC, B => WDIFF_3_net, C => 
        WDIFF_4_net, Y => OA1A_0_Y);
    
    AOI1_0 : AOI1
      port map(A => AND2_6_Y, B => NAND3A_1_Y, C => NOR3_0_Y, Y
         => AOI1_0_Y);
    
    AO1_10 : AO1
      port map(A => XOR2_35_Y, B => AND2_3_Y, C => AND2_1_Y, Y
         => AO1_10_Y);
    
    XOR2_35 : XOR2
      port map(A => MEM_WADDR_3_net, B => Fifo_rd_1_GND, Y => 
        XOR2_35_Y);
    
    DFN1P0_EMPTY : DFN1P0
      port map(D => EMPTYINT, CLK => PLL_Test1_0_Sys_66M_Clk, PRE
         => Main_ctl4SD_0_fifo_rst_n_3, Q => DFN1P0_EMPTY_0);
    
    AND2_17 : AND2
      port map(A => WBINNXTSHIFT_1_net, B => INV_3_Y, Y => 
        AND2_17_Y);
    
    DFN1E1C0_Q_40_inst : DFN1E1C0
      port map(D => QXI_40_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_2, E => DVLDI_1, Q => 
        \Z\\Fifo_rd_0_Q_[40]\\\);
    
    NOR2A_0 : NOR2A
      port map(A => MEM_RADDR_0_net, B => WBINNXTSHIFT_0_net, Y
         => NOR2A_0_Y);
    
    AO1_13 : AO1
      port map(A => XOR2_4_Y, B => AO1_8_Y, C => AND2_4_Y, Y => 
        AO1_13_Y);
    
    DFN1C0_MEM_WADDR_3_inst : DFN1C0
      port map(D => WBINNXTSHIFT_3_net, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => 
        Main_ctl4SD_0_fifo_rst_n_0, Q => MEM_WADDR_3_net);
    
    DFN1E1C0_Q_48_inst : DFN1E1C0
      port map(D => QXI_48_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_2, E => DVLDI_1, Q => 
        \Z\\Fifo_rd_0_Q_[48]\\\);
    
    DFN1E1C0_Q_9_inst : DFN1E1C0
      port map(D => QXI_9_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_3, E => DVLDI_2, Q => 
        \Z\\Fifo_rd_0_Q_[9]\\\);
    
    DFN1E1C0_Q_59_inst : DFN1E1C0
      port map(D => QXI_59_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_2, E => DVLDI_2, Q => 
        \Z\\Fifo_rd_0_Q_[59]\\\);
    
    XNOR2_WDIFF_1_inst : XNOR2
      port map(A => XOR2_14_Y, B => NOR2A_0_Y, Y => WDIFF_1_net);
    
    OR2A_0 : OR2A
      port map(A => Fifo_rd_1_GND, B => WDIFF_2_net, Y => 
        OR2A_0_Y);
    
    XNOR2_7 : XNOR2
      port map(A => MEM_RADDR_1_net, B => WBINNXTSHIFT_1_net, Y
         => XNOR2_7_Y);
    
    DFN1E1C0_Q_64_inst : DFN1E1C0
      port map(D => QXI_64_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_3, E => DVLDI_2, Q => 
        \Z\\Fifo_rd_0_Q_[64]\\\);
    
    DFN1C0_MEM_RADDR_2_inst : DFN1C0
      port map(D => RBINNXTSHIFT_2_net, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => 
        Main_ctl4SD_0_fifo_rst_n_0, Q => MEM_RADDR_2_net);
    
    AND2_4 : AND2
      port map(A => MEM_RADDR_2_net, B => Fifo_rd_1_GND, Y => 
        AND2_4_Y);
    
    AND2_FULLINT : AND2
      port map(A => AND2_7_Y, B => XOR2_23_Y, Y => FULLINT);
    
    DFN1C0_MEM_RADDR_1_inst : DFN1C0
      port map(D => RBINNXTSHIFT_1_net, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => 
        Main_ctl4SD_0_fifo_rst_n_0, Q => MEM_RADDR_1_net);
    
    XNOR2_5 : XNOR2
      port map(A => RBINNXTSHIFT_2_net, B => MEM_WADDR_2_net, Y
         => XNOR2_5_Y);
    
    DFN1E1C0_Q_21_inst : DFN1E1C0
      port map(D => QXI_21_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_1, E => DVLDI_0, Q => 
        \Z\\Fifo_rd_0_Q_[21]\\\);
    
    AO1_5 : AO1
      port map(A => AND2_24_Y, B => AO1_8_Y, C => AO1_11_Y, Y => 
        AO1_5_Y);
    
    DFN1E1C0_Q_50_inst : DFN1E1C0
      port map(D => QXI_50_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_2, E => DVLDI_1, Q => 
        \Z\\Fifo_rd_0_Q_[50]\\\);
    
    AND2_8 : AND2
      port map(A => MEM_WADDR_0_net, B => MEMORYWE, Y => AND2_8_Y);
    
    XOR2_3 : XOR2
      port map(A => WBINNXTSHIFT_3_net, B => INV_2_Y, Y => 
        XOR2_3_Y);
    
    RAM512X18_QXI_35_inst : RAM512X18
      port map(RADDR8 => Fifo_rd_1_GND, RADDR7 => Fifo_rd_1_GND, 
        RADDR6 => Fifo_rd_1_GND, RADDR5 => Fifo_rd_1_GND, RADDR4
         => Fifo_rd_1_GND, RADDR3 => MEM_RADDR_3_net, RADDR2 => 
        MEM_RADDR_2_net, RADDR1 => MEM_RADDR_1_net, RADDR0 => 
        MEM_RADDR_0_net, WADDR8 => Fifo_rd_1_GND, WADDR7 => 
        Fifo_rd_1_GND, WADDR6 => Fifo_rd_1_GND, WADDR5 => 
        Fifo_rd_1_GND, WADDR4 => Fifo_rd_1_GND, WADDR3 => 
        MEM_WADDR_3_net, WADDR2 => MEM_WADDR_2_net, WADDR1 => 
        MEM_WADDR_1_net, WADDR0 => MEM_WADDR_0_net, WD17 => 
        \Z\\Sdram_data_0_Sys_dataOut_[35]\\\, WD16 => 
        \Z\\Sdram_data_0_Sys_dataOut_[34]\\\, WD15 => 
        \Z\\Sdram_data_0_Sys_dataOut_[33]\\\, WD14 => 
        \Z\\Sdram_data_0_Sys_dataOut_[32]\\\, WD13 => 
        \Z\\Sdram_data_0_Sys_dataOut_[31]\\\, WD12 => 
        \Z\\Sdram_data_0_Sys_dataOut_[30]\\\, WD11 => 
        \Z\\Sdram_data_0_Sys_dataOut_[29]\\\, WD10 => 
        \Z\\Sdram_data_0_Sys_dataOut_[28]\\\, WD9 => 
        \Z\\Sdram_data_0_Sys_dataOut_[27]\\\, WD8 => 
        \Z\\Sdram_data_0_Sys_dataOut_[26]\\\, WD7 => 
        \Z\\Sdram_data_0_Sys_dataOut_[25]\\\, WD6 => 
        \Z\\Sdram_data_0_Sys_dataOut_[24]\\\, WD5 => 
        \Z\\Sdram_data_0_Sys_dataOut_[23]\\\, WD4 => 
        \Z\\Sdram_data_0_Sys_dataOut_[22]\\\, WD3 => 
        \Z\\Sdram_data_0_Sys_dataOut_[21]\\\, WD2 => 
        \Z\\Sdram_data_0_Sys_dataOut_[20]\\\, WD1 => 
        \Z\\Sdram_data_0_Sys_dataOut_[19]\\\, WD0 => 
        \Z\\Sdram_data_0_Sys_dataOut_[18]\\\, RW0 => 
        Fifo_rd_1_GND, RW1 => Fifo_rd_1_VCC, WW0 => Fifo_rd_1_GND, 
        WW1 => Fifo_rd_1_VCC, PIPE => Fifo_rd_1_GND, REN => 
        MEMRENEG, WEN => MEMWENEG, RCLK => 
        PLL_Test1_0_Sys_66M_Clk, WCLK => PLL_Test1_0_Sys_66M_Clk, 
        RESET => Main_ctl4SD_0_fifo_rst_n_3, RD17 => QXI_35_net, 
        RD16 => QXI_34_net, RD15 => QXI_33_net, RD14 => 
        QXI_32_net, RD13 => QXI_31_net, RD12 => QXI_30_net, RD11
         => QXI_29_net, RD10 => QXI_28_net, RD9 => QXI_27_net, 
        RD8 => QXI_26_net, RD7 => QXI_25_net, RD6 => QXI_24_net, 
        RD5 => QXI_23_net, RD4 => QXI_22_net, RD3 => QXI_21_net, 
        RD2 => QXI_20_net, RD1 => QXI_19_net, RD0 => QXI_18_net);
    
    DFN1E1C0_Q_31_inst : DFN1E1C0
      port map(D => QXI_31_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_1, E => DVLDI_1, Q => 
        \Z\\Fifo_rd_0_Q_[31]\\\);
    
    DFN1E1C0_Q_25_inst : DFN1E1C0
      port map(D => QXI_25_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_1, E => DVLDI_0, Q => 
        \Z\\Fifo_rd_0_Q_[25]\\\);
    
    DFN1E1C0_Q_58_inst : DFN1E1C0
      port map(D => QXI_58_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_2, E => DVLDI_2, Q => 
        \Z\\Fifo_rd_0_Q_[58]\\\);
    
    DFN1E1C0_Q_35_inst : DFN1E1C0
      port map(D => QXI_35_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_1, E => DVLDI_1, Q => 
        \Z\\Fifo_rd_0_Q_[35]\\\);
    
    DFN1E1C0_Q_19_inst : DFN1E1C0
      port map(D => QXI_19_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_1, E => DVLDI_0, Q => 
        \Z\\Fifo_rd_0_Q_[19]\\\);
    
    XOR2_28 : XOR2
      port map(A => MEM_RADDR_3_net, B => Fifo_rd_1_GND, Y => 
        XOR2_28_Y);
    
    XOR2_WDIFF_2_inst : XOR2
      port map(A => XOR2_20_Y, B => OR3_0_Y, Y => WDIFF_2_net);
    
    DFN1E1C0_Q_26_inst : DFN1E1C0
      port map(D => QXI_26_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_1, E => DVLDI_0, Q => 
        \Z\\Fifo_rd_0_Q_[26]\\\);
    
    DFN1E1C0_Q_22_inst : DFN1E1C0
      port map(D => QXI_22_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_1, E => DVLDI_0, Q => 
        \Z\\Fifo_rd_0_Q_[22]\\\);
    
    DFN1E1C0_Q_36_inst : DFN1E1C0
      port map(D => QXI_36_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_1, E => DVLDI_1, Q => 
        \Z\\Fifo_rd_0_Q_[36]\\\);
    
    AND2_21 : AND2
      port map(A => MEM_RADDR_3_net, B => Fifo_rd_1_GND, Y => 
        AND2_21_Y);
    
    XOR2_WDIFF_3_inst : XOR2
      port map(A => XOR2_9_Y, B => AO1_7_Y, Y => WDIFF_3_net);
    
    DFN1E1C0_Q_32_inst : DFN1E1C0
      port map(D => QXI_32_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_1, E => DVLDI_1, Q => 
        \Z\\Fifo_rd_0_Q_[32]\\\);
    
    DFN1E1C0_Q_6_inst : DFN1E1C0
      port map(D => QXI_6_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_3, E => DVLDI_2, Q => 
        \Z\\Fifo_rd_0_Q_[6]\\\);
    
    XOR2_0 : XOR2
      port map(A => MEM_WADDR_1_net, B => Fifo_rd_1_GND, Y => 
        XOR2_0_Y);
    
    NAND2_1 : NAND2
      port map(A => DFN1P0_EMPTY_0, B => Fifo_rd_1_VCC, Y => 
        NAND2_1_Y);
    
    DFN1E1C0_Q_44_inst : DFN1E1C0
      port map(D => QXI_44_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_2, E => DVLDI_1, Q => 
        \Z\\Fifo_rd_0_Q_[44]\\\);
    
    DFN1C0_MEM_RADDR_4_inst : DFN1C0
      port map(D => RBINNXTSHIFT_4_net, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => 
        Main_ctl4SD_0_fifo_rst_n_0, Q => MEM_RADDR_4_net);
    
    DFN1E1C0_Q_10_inst : DFN1E1C0
      port map(D => QXI_10_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_0, E => DVLDI_0, Q => 
        \Z\\Fifo_rd_0_Q_[10]\\\);
    
    AO1_4 : AO1
      port map(A => XOR2_11_Y, B => AO1_0_Y, C => AND2_3_Y, Y => 
        AO1_4_Y);
    
    DFN1E1C0_Q_71_inst : DFN1E1C0
      port map(D => QXI_71_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_3, E => DVLDI_2, Q => 
        \Z\\Fifo_rd_0_Q_[71]\\\);
    
    DFN1E1C0_Q_18_inst : DFN1E1C0
      port map(D => QXI_18_net, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => Main_ctl4SD_0_fifo_rst_n_0, E => DVLDI_0, Q => 
        \Z\\Fifo_rd_0_Q_[18]\\\);
    
    XOR2_36 : XOR2
      port map(A => MEM_RADDR_4_net, B => Fifo_rd_1_GND, Y => 
        XOR2_36_Y);
    
    XNOR2_8 : XNOR2
      port map(A => MEM_RADDR_3_net, B => WBINNXTSHIFT_3_net, Y
         => XNOR2_8_Y);
    
    XOR2_WDIFF_0_inst : XOR2
      port map(A => WBINNXTSHIFT_0_net, B => MEM_RADDR_0_net, Y
         => WDIFF_0_net);
    
    AND2_28 : AND2
      port map(A => MEM_RADDR_0_net, B => MEMORYRE, Y => 
        AND2_28_Y);
    
    AND2_25 : AND2
      port map(A => AND3_1_Y, B => XNOR2_6_Y, Y => AND2_25_Y);
    
    DFN1C0_DVLDI_RNI2T66_0 : BUFF
      port map(A => DVLDI, Y => DVLDI_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3;
use proasic3.all;

entity Sdram_data is

    port( Sd_DQ_in                             : in    std_logic_vector(71 downto 0);
          \Z\\Sdram_data_0_Sys_dataOut_[71]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[70]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[69]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[68]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[67]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[66]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[65]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[64]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[63]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[62]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[61]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[60]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[59]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[58]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[57]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[56]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[55]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[54]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[53]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[52]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[51]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[50]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[49]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[48]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[47]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[46]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[45]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[44]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[43]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[42]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[41]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[40]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[39]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[38]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[37]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[36]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[35]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[34]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[33]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[32]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[31]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[30]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[29]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[28]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[27]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[26]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[25]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[24]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[23]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[22]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[21]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[20]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[19]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[18]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[17]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[16]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[15]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[14]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[13]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[12]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[11]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[10]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[9]\\\  : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[8]\\\  : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[7]\\\  : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[6]\\\  : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[5]\\\  : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[4]\\\  : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[3]\\\  : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[2]\\\  : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[1]\\\  : out   std_logic;
          PLL_Test1_0_SysRst_O                 : in    std_logic;
          PLL_Test1_0_Sys_66M_Clk              : in    std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[0]\\\  : out   std_logic;
          \Z\\SDram_rd_0_rd_state_[1]\\\       : in    std_logic;
          \Z\\SDram_rd_0_rd_state_[2]\\\       : in    std_logic;
          \Z\\SDram_rd_0_rd_state_[0]\\\       : in    std_logic
        );

end Sdram_data;

architecture DEF_ARCH of Sdram_data is 

  component DFN1E1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal \sys_dataout5_1\, \sys_dataout5_0\, \sys_dataout5\, 
        \GND\, \VCC\, GND_0, VCC_0 : std_logic;

begin 


    \Sys_dataOut[25]\ : DFN1E1C0
      port map(D => Sd_DQ_in(25), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5_0\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[25]\\\);
    
    \Sys_dataOut[54]\ : DFN1E1C0
      port map(D => Sd_DQ_in(54), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[54]\\\);
    
    \Sys_dataOut[29]\ : DFN1E1C0
      port map(D => Sd_DQ_in(29), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5_0\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[29]\\\);
    
    \Sys_dataOut[36]\ : DFN1E1C0
      port map(D => Sd_DQ_in(36), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5_1\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[36]\\\);
    
    \Sys_dataOut[64]\ : DFN1E1C0
      port map(D => Sd_DQ_in(64), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[64]\\\);
    
    \Sys_dataOut[3]\ : DFN1E1C0
      port map(D => Sd_DQ_in(3), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5_1\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[3]\\\);
    
    sys_dataout5_1 : NOR3B
      port map(A => \Z\\SDram_rd_0_rd_state_[0]\\\, B => 
        \Z\\SDram_rd_0_rd_state_[2]\\\, C => 
        \Z\\SDram_rd_0_rd_state_[1]\\\, Y => \sys_dataout5_1\);
    
    \Sys_dataOut[46]\ : DFN1E1C0
      port map(D => Sd_DQ_in(46), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5_1\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[46]\\\);
    
    \Sys_dataOut[30]\ : DFN1E1C0
      port map(D => Sd_DQ_in(30), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5_0\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[30]\\\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \Sys_dataOut[37]\ : DFN1E1C0
      port map(D => Sd_DQ_in(37), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5_1\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[37]\\\);
    
    \Sys_dataOut[18]\ : DFN1E1C0
      port map(D => Sd_DQ_in(18), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5_0\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[18]\\\);
    
    \Sys_dataOut[40]\ : DFN1E1C0
      port map(D => Sd_DQ_in(40), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5_1\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[40]\\\);
    
    \Sys_dataOut[11]\ : DFN1E1C0
      port map(D => Sd_DQ_in(11), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5_0\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[11]\\\);
    
    \Sys_dataOut[12]\ : DFN1E1C0
      port map(D => Sd_DQ_in(12), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5_0\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[12]\\\);
    
    \Sys_dataOut[47]\ : DFN1E1C0
      port map(D => Sd_DQ_in(47), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5_1\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[47]\\\);
    
    \Sys_dataOut[35]\ : DFN1E1C0
      port map(D => Sd_DQ_in(35), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5_1\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[35]\\\);
    
    \Sys_dataOut[56]\ : DFN1E1C0
      port map(D => Sd_DQ_in(56), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[56]\\\);
    
    \Sys_dataOut[66]\ : DFN1E1C0
      port map(D => Sd_DQ_in(66), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[66]\\\);
    
    \Sys_dataOut[39]\ : DFN1E1C0
      port map(D => Sd_DQ_in(39), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5_1\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[39]\\\);
    
    \Sys_dataOut[45]\ : DFN1E1C0
      port map(D => Sd_DQ_in(45), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5_1\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[45]\\\);
    
    \Sys_dataOut[5]\ : DFN1E1C0
      port map(D => Sd_DQ_in(5), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[5]\\\);
    
    \Sys_dataOut[50]\ : DFN1E1C0
      port map(D => Sd_DQ_in(50), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5_1\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[50]\\\);
    
    \Sys_dataOut[71]\ : DFN1E1C0
      port map(D => Sd_DQ_in(71), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[71]\\\);
    
    \Sys_dataOut[13]\ : DFN1E1C0
      port map(D => Sd_DQ_in(13), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5_0\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[13]\\\);
    
    \Sys_dataOut[57]\ : DFN1E1C0
      port map(D => Sd_DQ_in(57), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[57]\\\);
    
    \Sys_dataOut[49]\ : DFN1E1C0
      port map(D => Sd_DQ_in(49), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5_1\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[49]\\\);
    
    \Sys_dataOut[28]\ : DFN1E1C0
      port map(D => Sd_DQ_in(28), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5_0\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[28]\\\);
    
    \Sys_dataOut[60]\ : DFN1E1C0
      port map(D => Sd_DQ_in(60), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[60]\\\);
    
    \Sys_dataOut[21]\ : DFN1E1C0
      port map(D => Sd_DQ_in(21), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5_0\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[21]\\\);
    
    \Sys_dataOut[67]\ : DFN1E1C0
      port map(D => Sd_DQ_in(67), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[67]\\\);
    
    \Sys_dataOut[22]\ : DFN1E1C0
      port map(D => Sd_DQ_in(22), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5_0\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[22]\\\);
    
    \Sys_dataOut[55]\ : DFN1E1C0
      port map(D => Sd_DQ_in(55), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[55]\\\);
    
    \Sys_dataOut[65]\ : DFN1E1C0
      port map(D => Sd_DQ_in(65), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[65]\\\);
    
    \Sys_dataOut[8]\ : DFN1E1C0
      port map(D => Sd_DQ_in(8), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[8]\\\);
    
    \Sys_dataOut[59]\ : DFN1E1C0
      port map(D => Sd_DQ_in(59), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[59]\\\);
    
    \Sys_dataOut[1]\ : DFN1E1C0
      port map(D => Sd_DQ_in(1), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5_0\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[1]\\\);
    
    \Sys_dataOut[14]\ : DFN1E1C0
      port map(D => Sd_DQ_in(14), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5_0\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[14]\\\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \Sys_dataOut[69]\ : DFN1E1C0
      port map(D => Sd_DQ_in(69), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[69]\\\);
    
    \Sys_dataOut[23]\ : DFN1E1C0
      port map(D => Sd_DQ_in(23), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5_0\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[23]\\\);
    
    \Sys_dataOut[0]\ : DFN1E1C0
      port map(D => Sd_DQ_in(0), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5_0\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[0]\\\);
    
    sys_dataout5_0 : NOR3B
      port map(A => \Z\\SDram_rd_0_rd_state_[0]\\\, B => 
        \Z\\SDram_rd_0_rd_state_[2]\\\, C => 
        \Z\\SDram_rd_0_rd_state_[1]\\\, Y => \sys_dataout5_0\);
    
    \Sys_dataOut[2]\ : DFN1E1C0
      port map(D => Sd_DQ_in(2), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5_0\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[2]\\\);
    
    \Sys_dataOut[38]\ : DFN1E1C0
      port map(D => Sd_DQ_in(38), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5_1\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[38]\\\);
    
    \Sys_dataOut[31]\ : DFN1E1C0
      port map(D => Sd_DQ_in(31), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5_1\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[31]\\\);
    
    \Sys_dataOut[32]\ : DFN1E1C0
      port map(D => Sd_DQ_in(32), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5_1\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[32]\\\);
    
    \Sys_dataOut[4]\ : DFN1E1C0
      port map(D => Sd_DQ_in(4), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5_1\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[4]\\\);
    
    \Sys_dataOut[9]\ : DFN1E1C0
      port map(D => Sd_DQ_in(9), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[9]\\\);
    
    \Sys_dataOut[6]\ : DFN1E1C0
      port map(D => Sd_DQ_in(6), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[6]\\\);
    
    \Sys_dataOut[48]\ : DFN1E1C0
      port map(D => Sd_DQ_in(48), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5_1\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[48]\\\);
    
    \Sys_dataOut[24]\ : DFN1E1C0
      port map(D => Sd_DQ_in(24), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5_0\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[24]\\\);
    
    sys_dataout5 : NOR3B
      port map(A => \Z\\SDram_rd_0_rd_state_[0]\\\, B => 
        \Z\\SDram_rd_0_rd_state_[2]\\\, C => 
        \Z\\SDram_rd_0_rd_state_[1]\\\, Y => \sys_dataout5\);
    
    \Sys_dataOut[41]\ : DFN1E1C0
      port map(D => Sd_DQ_in(41), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5_1\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[41]\\\);
    
    \Sys_dataOut[42]\ : DFN1E1C0
      port map(D => Sd_DQ_in(42), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5_1\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[42]\\\);
    
    \Sys_dataOut[16]\ : DFN1E1C0
      port map(D => Sd_DQ_in(16), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5_0\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[16]\\\);
    
    \Sys_dataOut[7]\ : DFN1E1C0
      port map(D => Sd_DQ_in(7), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[7]\\\);
    
    \Sys_dataOut[33]\ : DFN1E1C0
      port map(D => Sd_DQ_in(33), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5_1\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[33]\\\);
    
    \Sys_dataOut[58]\ : DFN1E1C0
      port map(D => Sd_DQ_in(58), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[58]\\\);
    
    \Sys_dataOut[10]\ : DFN1E1C0
      port map(D => Sd_DQ_in(10), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5_0\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[10]\\\);
    
    \Sys_dataOut[51]\ : DFN1E1C0
      port map(D => Sd_DQ_in(51), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5_1\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[51]\\\);
    
    \Sys_dataOut[17]\ : DFN1E1C0
      port map(D => Sd_DQ_in(17), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5_0\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[17]\\\);
    
    \Sys_dataOut[68]\ : DFN1E1C0
      port map(D => Sd_DQ_in(68), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[68]\\\);
    
    \Sys_dataOut[52]\ : DFN1E1C0
      port map(D => Sd_DQ_in(52), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5_1\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[52]\\\);
    
    \Sys_dataOut[43]\ : DFN1E1C0
      port map(D => Sd_DQ_in(43), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5_1\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[43]\\\);
    
    \Sys_dataOut[61]\ : DFN1E1C0
      port map(D => Sd_DQ_in(61), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[61]\\\);
    
    \Sys_dataOut[62]\ : DFN1E1C0
      port map(D => Sd_DQ_in(62), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[62]\\\);
    
    \Sys_dataOut[26]\ : DFN1E1C0
      port map(D => Sd_DQ_in(26), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5_0\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[26]\\\);
    
    \Sys_dataOut[15]\ : DFN1E1C0
      port map(D => Sd_DQ_in(15), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5_0\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[15]\\\);
    
    \Sys_dataOut[70]\ : DFN1E1C0
      port map(D => Sd_DQ_in(70), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[70]\\\);
    
    \Sys_dataOut[34]\ : DFN1E1C0
      port map(D => Sd_DQ_in(34), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5_1\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[34]\\\);
    
    \Sys_dataOut[19]\ : DFN1E1C0
      port map(D => Sd_DQ_in(19), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5_0\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[19]\\\);
    
    \Sys_dataOut[53]\ : DFN1E1C0
      port map(D => Sd_DQ_in(53), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[53]\\\);
    
    \Sys_dataOut[20]\ : DFN1E1C0
      port map(D => Sd_DQ_in(20), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5_0\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[20]\\\);
    
    \Sys_dataOut[44]\ : DFN1E1C0
      port map(D => Sd_DQ_in(44), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5_1\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[44]\\\);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    \Sys_dataOut[63]\ : DFN1E1C0
      port map(D => Sd_DQ_in(63), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[63]\\\);
    
    \Sys_dataOut[27]\ : DFN1E1C0
      port map(D => Sd_DQ_in(27), CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, E => \sys_dataout5_0\, Q => 
        \Z\\Sdram_data_0_Sys_dataOut_[27]\\\);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3;
use proasic3.all;

entity adc_muxtmp_test is

    port( PLL_Test1_0_SysRst_O                        : in    std_logic;
          PLL_Test1_0_Sys_66M_Clk                     : in    std_logic;
          CMOS_DrvX_0_AdcEn                           : in    std_logic;
          \Z\\adc_muxtmp_test_0_DataOut41to28_[29]\\\ : out   std_logic;
          \Z\\adc_muxtmp_test_0_DataOut27to14_[14]\\\ : out   std_logic;
          \Z\\adc_muxtmp_test_0_DataOut55to42_[43]\\\ : out   std_logic
        );

end adc_muxtmp_test;

architecture DEF_ARCH of adc_muxtmp_test is 

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AO1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XA1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component AO1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \DataOut_1_RNO[42]_net_1\, \ChSel[1]_net_1\, 
        \ChSel[0]_net_1\, \DataOut_1_RNO[14]_net_1\, 
        \DataOut_1_RNO[29]_net_1\, \ChSel_3[0]\, \ChSel_3[1]\, 
        \Z\\adc_muxtmp_test_0_DataOut41to28_[29]\\_net_1\, 
        \Z\\adc_muxtmp_test_0_DataOut27to14_[14]\\_net_1\, 
        \Z\\adc_muxtmp_test_0_DataOut55to42_[43]\\_net_1\, \GND\, 
        \VCC\, GND_0, VCC_0 : std_logic;

begin 

    \Z\\adc_muxtmp_test_0_DataOut41to28_[29]\\\ <= 
        \Z\\adc_muxtmp_test_0_DataOut41to28_[29]\\_net_1\;
    \Z\\adc_muxtmp_test_0_DataOut27to14_[14]\\\ <= 
        \Z\\adc_muxtmp_test_0_DataOut27to14_[14]\\_net_1\;
    \Z\\adc_muxtmp_test_0_DataOut55to42_[43]\\\ <= 
        \Z\\adc_muxtmp_test_0_DataOut55to42_[43]\\_net_1\;

    \ChSel[0]\ : DFN1C0
      port map(D => \ChSel_3[0]\, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \ChSel[0]_net_1\);
    
    \DataOut_1_RNO[14]\ : AO1A
      port map(A => \ChSel[1]_net_1\, B => \ChSel[0]_net_1\, C
         => \Z\\adc_muxtmp_test_0_DataOut27to14_[14]\\_net_1\, Y
         => \DataOut_1_RNO[14]_net_1\);
    
    \ChSel_RNO[1]\ : XA1B
      port map(A => \ChSel[0]_net_1\, B => \ChSel[1]_net_1\, C
         => CMOS_DrvX_0_AdcEn, Y => \ChSel_3[1]\);
    
    \DataOut_1[29]\ : DFN1C0
      port map(D => \DataOut_1_RNO[29]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \Z\\adc_muxtmp_test_0_DataOut41to28_[29]\\_net_1\);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    \ChSel_RNO[0]\ : NOR2
      port map(A => \ChSel[0]_net_1\, B => CMOS_DrvX_0_AdcEn, Y
         => \ChSel_3[0]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \DataOut_1_RNO[29]\ : AO1A
      port map(A => \ChSel[0]_net_1\, B => \ChSel[1]_net_1\, C
         => \Z\\adc_muxtmp_test_0_DataOut41to28_[29]\\_net_1\, Y
         => \DataOut_1_RNO[29]_net_1\);
    
    \DataOut_1[42]\ : DFN1C0
      port map(D => \DataOut_1_RNO[42]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \Z\\adc_muxtmp_test_0_DataOut55to42_[43]\\_net_1\);
    
    \DataOut_1[14]\ : DFN1C0
      port map(D => \DataOut_1_RNO[14]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \Z\\adc_muxtmp_test_0_DataOut27to14_[14]\\_net_1\);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \DataOut_1_RNO[42]\ : AO1
      port map(A => \ChSel[1]_net_1\, B => \ChSel[0]_net_1\, C
         => \Z\\adc_muxtmp_test_0_DataOut55to42_[43]\\_net_1\, Y
         => \DataOut_1_RNO[42]_net_1\);
    
    \ChSel[1]\ : DFN1C0
      port map(D => \ChSel_3[1]\, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \ChSel[1]_net_1\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3;
use proasic3.all;

entity my_pll is

    port( my_pll_VCC              : in    std_logic;
          my_pll_GND              : in    std_logic;
          ExterCLk_c              : in    std_logic;
          PLL_Lock                : out   std_logic;
          PLL_Test1_0_Sdram_clk   : out   std_logic;
          PLL_Test1_0_ADC_66M_Clk : out   std_logic;
          PLL_Test1_0_Sys_66M_Clk : out   std_logic
        );

end my_pll;

architecture DEF_ARCH of my_pll is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component PLL
    generic (VCOFREQUENCY:real := 0.0);

    port( CLKA      : in    std_logic := 'U';
          EXTFB     : in    std_logic := 'U';
          POWERDOWN : in    std_logic := 'U';
          GLA       : out   std_logic;
          LOCK      : out   std_logic;
          GLB       : out   std_logic;
          YB        : out   std_logic;
          GLC       : out   std_logic;
          YC        : out   std_logic;
          OADIV0    : in    std_logic := 'U';
          OADIV1    : in    std_logic := 'U';
          OADIV2    : in    std_logic := 'U';
          OADIV3    : in    std_logic := 'U';
          OADIV4    : in    std_logic := 'U';
          OAMUX0    : in    std_logic := 'U';
          OAMUX1    : in    std_logic := 'U';
          OAMUX2    : in    std_logic := 'U';
          DLYGLA0   : in    std_logic := 'U';
          DLYGLA1   : in    std_logic := 'U';
          DLYGLA2   : in    std_logic := 'U';
          DLYGLA3   : in    std_logic := 'U';
          DLYGLA4   : in    std_logic := 'U';
          OBDIV0    : in    std_logic := 'U';
          OBDIV1    : in    std_logic := 'U';
          OBDIV2    : in    std_logic := 'U';
          OBDIV3    : in    std_logic := 'U';
          OBDIV4    : in    std_logic := 'U';
          OBMUX0    : in    std_logic := 'U';
          OBMUX1    : in    std_logic := 'U';
          OBMUX2    : in    std_logic := 'U';
          DLYYB0    : in    std_logic := 'U';
          DLYYB1    : in    std_logic := 'U';
          DLYYB2    : in    std_logic := 'U';
          DLYYB3    : in    std_logic := 'U';
          DLYYB4    : in    std_logic := 'U';
          DLYGLB0   : in    std_logic := 'U';
          DLYGLB1   : in    std_logic := 'U';
          DLYGLB2   : in    std_logic := 'U';
          DLYGLB3   : in    std_logic := 'U';
          DLYGLB4   : in    std_logic := 'U';
          OCDIV0    : in    std_logic := 'U';
          OCDIV1    : in    std_logic := 'U';
          OCDIV2    : in    std_logic := 'U';
          OCDIV3    : in    std_logic := 'U';
          OCDIV4    : in    std_logic := 'U';
          OCMUX0    : in    std_logic := 'U';
          OCMUX1    : in    std_logic := 'U';
          OCMUX2    : in    std_logic := 'U';
          DLYYC0    : in    std_logic := 'U';
          DLYYC1    : in    std_logic := 'U';
          DLYYC2    : in    std_logic := 'U';
          DLYYC3    : in    std_logic := 'U';
          DLYYC4    : in    std_logic := 'U';
          DLYGLC0   : in    std_logic := 'U';
          DLYGLC1   : in    std_logic := 'U';
          DLYGLC2   : in    std_logic := 'U';
          DLYGLC3   : in    std_logic := 'U';
          DLYGLC4   : in    std_logic := 'U';
          FINDIV0   : in    std_logic := 'U';
          FINDIV1   : in    std_logic := 'U';
          FINDIV2   : in    std_logic := 'U';
          FINDIV3   : in    std_logic := 'U';
          FINDIV4   : in    std_logic := 'U';
          FINDIV5   : in    std_logic := 'U';
          FINDIV6   : in    std_logic := 'U';
          FBDIV0    : in    std_logic := 'U';
          FBDIV1    : in    std_logic := 'U';
          FBDIV2    : in    std_logic := 'U';
          FBDIV3    : in    std_logic := 'U';
          FBDIV4    : in    std_logic := 'U';
          FBDIV5    : in    std_logic := 'U';
          FBDIV6    : in    std_logic := 'U';
          FBDLY0    : in    std_logic := 'U';
          FBDLY1    : in    std_logic := 'U';
          FBDLY2    : in    std_logic := 'U';
          FBDLY3    : in    std_logic := 'U';
          FBDLY4    : in    std_logic := 'U';
          FBSEL0    : in    std_logic := 'U';
          FBSEL1    : in    std_logic := 'U';
          XDLYSEL   : in    std_logic := 'U';
          VCOSEL0   : in    std_logic := 'U';
          VCOSEL1   : in    std_logic := 'U';
          VCOSEL2   : in    std_logic := 'U'
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

    signal Core_YB, Core_YC, \GND\, \VCC\, GND_0, VCC_0
         : std_logic;

begin 


    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    Core : PLL
      generic map(VCOFREQUENCY => 66.0)

      port map(CLKA => ExterCLk_c, EXTFB => my_pll_GND, POWERDOWN
         => my_pll_VCC, GLA => PLL_Test1_0_Sys_66M_Clk, LOCK => 
        PLL_Lock, GLB => PLL_Test1_0_ADC_66M_Clk, YB => Core_YB, 
        GLC => PLL_Test1_0_Sdram_clk, YC => Core_YC, OADIV0 => 
        my_pll_GND, OADIV1 => my_pll_GND, OADIV2 => my_pll_GND, 
        OADIV3 => my_pll_GND, OADIV4 => my_pll_GND, OAMUX0 => 
        my_pll_GND, OAMUX1 => my_pll_GND, OAMUX2 => my_pll_VCC, 
        DLYGLA0 => my_pll_GND, DLYGLA1 => my_pll_GND, DLYGLA2 => 
        my_pll_GND, DLYGLA3 => my_pll_GND, DLYGLA4 => my_pll_GND, 
        OBDIV0 => my_pll_GND, OBDIV1 => my_pll_GND, OBDIV2 => 
        my_pll_GND, OBDIV3 => my_pll_GND, OBDIV4 => my_pll_GND, 
        OBMUX0 => my_pll_VCC, OBMUX1 => my_pll_GND, OBMUX2 => 
        my_pll_VCC, DLYYB0 => my_pll_GND, DLYYB1 => my_pll_GND, 
        DLYYB2 => my_pll_GND, DLYYB3 => my_pll_GND, DLYYB4 => 
        my_pll_GND, DLYGLB0 => my_pll_GND, DLYGLB1 => my_pll_GND, 
        DLYGLB2 => my_pll_VCC, DLYGLB3 => my_pll_GND, DLYGLB4 => 
        my_pll_GND, OCDIV0 => my_pll_GND, OCDIV1 => my_pll_GND, 
        OCDIV2 => my_pll_GND, OCDIV3 => my_pll_GND, OCDIV4 => 
        my_pll_GND, OCMUX0 => my_pll_GND, OCMUX1 => my_pll_VCC, 
        OCMUX2 => my_pll_GND, DLYYC0 => my_pll_GND, DLYYC1 => 
        my_pll_GND, DLYYC2 => my_pll_GND, DLYYC3 => my_pll_GND, 
        DLYYC4 => my_pll_GND, DLYGLC0 => my_pll_GND, DLYGLC1 => 
        my_pll_GND, DLYGLC2 => my_pll_GND, DLYGLC3 => my_pll_VCC, 
        DLYGLC4 => my_pll_GND, FINDIV0 => my_pll_VCC, FINDIV1 => 
        my_pll_VCC, FINDIV2 => my_pll_GND, FINDIV3 => my_pll_VCC, 
        FINDIV4 => my_pll_GND, FINDIV5 => my_pll_GND, FINDIV6 => 
        my_pll_GND, FBDIV0 => my_pll_VCC, FBDIV1 => my_pll_VCC, 
        FBDIV2 => my_pll_GND, FBDIV3 => my_pll_VCC, FBDIV4 => 
        my_pll_GND, FBDIV5 => my_pll_GND, FBDIV6 => my_pll_GND, 
        FBDLY0 => my_pll_GND, FBDLY1 => my_pll_GND, FBDLY2 => 
        my_pll_GND, FBDLY3 => my_pll_GND, FBDLY4 => my_pll_GND, 
        FBSEL0 => my_pll_VCC, FBSEL1 => my_pll_GND, XDLYSEL => 
        my_pll_GND, VCOSEL0 => my_pll_VCC, VCOSEL1 => my_pll_VCC, 
        VCOSEL2 => my_pll_GND);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3;
use proasic3.all;

entity PLL_Test1 is

    port( PLL_Test1_0_ADC_66M_Clk : out   std_logic;
          PLL_Test1_0_Sdram_clk   : out   std_logic;
          ExterCLk_c              : in    std_logic;
          PLL_Test1_GND           : in    std_logic;
          PLL_Test1_0_SysRst_O    : out   std_logic;
          PLL_Test1_VCC           : in    std_logic;
          PLL_Test1_0_Sys_66M_Clk : out   std_logic
        );

end PLL_Test1;

architecture DEF_ARCH of PLL_Test1 is 

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component my_pll
    port( my_pll_VCC              : in    std_logic := 'U';
          my_pll_GND              : in    std_logic := 'U';
          ExterCLk_c              : in    std_logic := 'U';
          PLL_Lock                : out   std_logic;
          PLL_Test1_0_Sdram_clk   : out   std_logic;
          PLL_Test1_0_ADC_66M_Clk : out   std_logic;
          PLL_Test1_0_Sys_66M_Clk : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component CLKINT
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \RstBuf[0]_net_1\, PLL_Lock, \RstBuf[1]_net_1\, 
        \PLL_Test1_0_Sys_66M_Clk\, \GND\, \VCC\, GND_0, VCC_0
         : std_logic;

    for all : my_pll
	Use entity work.my_pll(DEF_ARCH);
begin 

    PLL_Test1_0_Sys_66M_Clk <= \PLL_Test1_0_Sys_66M_Clk\;

    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    Module_my_pll : my_pll
      port map(my_pll_VCC => PLL_Test1_VCC, my_pll_GND => 
        PLL_Test1_GND, ExterCLk_c => ExterCLk_c, PLL_Lock => 
        PLL_Lock, PLL_Test1_0_Sdram_clk => PLL_Test1_0_Sdram_clk, 
        PLL_Test1_0_ADC_66M_Clk => PLL_Test1_0_ADC_66M_Clk, 
        PLL_Test1_0_Sys_66M_Clk => \PLL_Test1_0_Sys_66M_Clk\);
    
    \RstBuf[0]\ : DFN1C0
      port map(D => PLL_Test1_VCC, CLK => 
        \PLL_Test1_0_Sys_66M_Clk\, CLR => PLL_Lock, Q => 
        \RstBuf[0]_net_1\);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    Module_CLKINT : CLKINT
      port map(A => \RstBuf[1]_net_1\, Y => PLL_Test1_0_SysRst_O);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \RstBuf[1]\ : DFN1C0
      port map(D => \RstBuf[0]_net_1\, CLK => 
        \PLL_Test1_0_Sys_66M_Clk\, CLR => PLL_Lock, Q => 
        \RstBuf[1]_net_1\);
    
    GND_i : GND
      port map(Y => \GND\);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3;
use proasic3.all;

entity Sdram_ctl_v2 is

    port( SD_cke_c_c                   : out   std_logic_vector(0 to 0);
          pr_state_ns_3                : out   std_logic;
          Sdram_ini_0_Sd_iniOK_i       : in    std_logic;
          Sdram_ctl_v2_0_SD_iniEn      : out   std_logic;
          Sdram_ctl_v2_0_SD_RefEn      : out   std_logic;
          Sdram_ctl_v2_0_SD_rdEN_noact : out   std_logic;
          PLL_Test1_0_SysRst_O         : in    std_logic;
          PLL_Test1_0_Sys_66M_Clk      : in    std_logic;
          Sdram_ctl_v2_0_SD_pdEN       : out   std_logic;
          Fifo_wr_0_AFULL              : in    std_logic;
          SDRAM_wr_0_SD_WrOK           : in    std_logic;
          ref_ok_2                     : in    std_logic;
          ref_ok_1                     : in    std_logic;
          CMOS_DrvX_0_LVDSen_2         : in    std_logic;
          CMOS_DrvX_0_SDramEn_0        : in    std_logic;
          Sdram_ini_0_Sd_iniOK         : in    std_logic;
          Fifo_rd_0_AFULL              : in    std_logic;
          CMOS_DrvX_0_LVDSen_1         : in    std_logic;
          SDram_rd_0_SD_RdOK           : in    std_logic;
          Sdram_ctl_v2_0_SD_rdEn       : out   std_logic;
          Sdram_ctl_v2_0_SD_rdEn_i     : out   std_logic;
          Sdram_ctl_v2_0_SD_wrEn       : out   std_logic;
          Sdram_ctl_v2_0_SD_wrEn_i     : out   std_logic
        );

end Sdram_ctl_v2;

architecture DEF_ARCH of Sdram_ctl_v2 is 

  component XNOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component OAI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OA1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1E0C0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          CLR : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component AOI1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component OR3A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AOI1B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component INV
    port( A : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component AX1C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component DFN1P0
    port( D   : in    std_logic := 'U';
          CLK : in    std_logic := 'U';
          PRE : in    std_logic := 'U';
          Q   : out   std_logic
        );
  end component;

  component MX2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          S : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR3C
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component AO1A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3B
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component NOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component OR2A
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal \pr_state_ns_i[8]\, \pr_state_ns_i_0[3]\, 
        \pr_state_RNITULC[11]_net_1\, N_164, N_177, un2lto11_0, 
        \temp[10]_net_1\, \temp[11]_net_1\, 
        \pr_state_ns_i_a2_0[7]\, \pr_state[4]_net_1\, 
        \pr_state[7]_net_1\, un2lto9_0, \temp[8]_net_1\, 
        \temp[9]_net_1\, un2lto7_1, \temp[6]_net_1\, 
        \temp[5]_net_1\, \temp[7]_net_1\, un2lto4_0, 
        \temp[3]_net_1\, \temp[4]_net_1\, un2, un2lt9, un2lt4, 
        N_169, \pr_state[11]_net_1\, \pr_state[0]_net_1\, N_162, 
        N_171, \pr_state[6]_net_1\, N_172, \pr_state[10]_net_1\, 
        \pr_state[5]_net_1\, N_163, N_173, \pr_state[9]_net_1\, 
        N_178, \pr_state[8]_net_1\, N_182, N_160, 
        \pr_state_RNO[9]_net_1\, \pr_state_ns[8]\, N_174, N_175, 
        \pr_state_RNO_0[2]\, \pr_state_ns[6]\, \pr_state_ns_2[6]\, 
        \pr_state_RNO[8]_net_1\, \pr_state_RNO[4]_net_1\, 
        \pr_state_ns_i_0[7]\, \pr_state_RNO[10]_net_1\, 
        \pr_state_RNO[11]_net_1\, \pr_state_ns_i_a2_1_0[7]\, 
        \pr_state_ns_i_a2_0_0[7]\, \temp_10\, temp_n10, 
        \PowerOK_RNO\, \temp_c2\, \temp[0]_net_1\, 
        \temp[1]_net_1\, \temp[2]_net_1\, \temp_c4\, \temp_c8\, 
        \temp_c6\, \temp_c9\, temp_n1, temp_n2, temp_n3, temp_n4, 
        temp_n5, temp_n7, temp_n8, temp_n9, \temp_20_0\, temp_n11, 
        temp_n6, \pr_state_ns[5]\, N_159, N_167, 
        \pr_state_RNO[0]_net_1\, \pr_state[1]_net_1\, 
        \pr_state_RNO_0[1]\, \pr_state[2]_net_1\, 
        \pr_state_RNO[7]_net_1\, \pr_state[3]_net_1\, 
        \SD_RefEn_RNO\, SD_iniEn_1_sqmuxa, \SD_cke_c_c[0]\, 
        \Sdram_ctl_v2_0_SD_wrEn\, \Sdram_ctl_v2_0_SD_rdEn\, \GND\, 
        \VCC\, GND_0, VCC_0 : std_logic;

begin 

    SD_cke_c_c(0) <= \SD_cke_c_c[0]\;
    pr_state_ns_3 <= \pr_state_ns[8]\;
    Sdram_ctl_v2_0_SD_rdEn <= \Sdram_ctl_v2_0_SD_rdEn\;
    Sdram_ctl_v2_0_SD_wrEn <= \Sdram_ctl_v2_0_SD_wrEn\;

    temp_n3_0 : XNOR2
      port map(A => \temp_c2\, B => \temp[3]_net_1\, Y => temp_n3);
    
    \pr_state_RNO[11]\ : NOR3A
      port map(A => \pr_state_ns[8]\, B => N_169, C => N_171, Y
         => \pr_state_RNO[11]_net_1\);
    
    \pr_state_RNO_0[9]\ : OA1C
      port map(A => \pr_state[9]_net_1\, B => SDRAM_wr_0_SD_WrOK, 
        C => \pr_state[6]_net_1\, Y => N_174);
    
    \pr_state[11]\ : DFN1C0
      port map(D => \pr_state_RNO[11]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \pr_state[11]_net_1\);
    
    \pr_state_RNIQKC1[8]\ : OAI1
      port map(A => ref_ok_1, B => ref_ok_2, C => 
        \pr_state[8]_net_1\, Y => N_160);
    
    \temp_RNISK0M1[10]\ : OA1
      port map(A => un2lt9, B => un2lto9_0, C => un2lto11_0, Y
         => un2);
    
    \temp_RNI1OEF[6]\ : NOR3C
      port map(A => \temp[6]_net_1\, B => \temp[5]_net_1\, C => 
        \temp[7]_net_1\, Y => un2lto7_1);
    
    SD_iniEn_RNO : NOR2
      port map(A => Sdram_ini_0_Sd_iniOK, B => \SD_cke_c_c[0]\, Y
         => SD_iniEn_1_sqmuxa);
    
    SD_iniEn : DFN1E0C0
      port map(D => Sdram_ini_0_Sd_iniOK_i, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, E
         => SD_iniEn_1_sqmuxa, Q => Sdram_ctl_v2_0_SD_iniEn);
    
    \pr_state_RNO_0[4]\ : OA1C
      port map(A => CMOS_DrvX_0_LVDSen_1, B => N_160, C => 
        \pr_state_ns_i_a2_0[7]\, Y => N_182);
    
    SD_wrEn : DFN1C0
      port map(D => \pr_state[9]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \Sdram_ctl_v2_0_SD_wrEn\);
    
    SD_rdEN_noact : DFN1C0
      port map(D => \pr_state[10]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => Sdram_ctl_v2_0_SD_rdEN_noact);
    
    \temp[9]\ : DFN1E0C0
      port map(D => temp_n9, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => un2, Q => \temp[9]_net_1\);
    
    \pr_state_RNO_1[4]\ : AOI1
      port map(A => \pr_state_ns_i_a2_1_0[7]\, B => 
        \pr_state_ns_i_a2_0_0[7]\, C => \pr_state[8]_net_1\, Y
         => \pr_state_ns_i_0[7]\);
    
    \temp_RNITBH2[10]\ : NOR2B
      port map(A => \temp[10]_net_1\, B => \temp[11]_net_1\, Y
         => un2lto11_0);
    
    temp_n8_0 : AX1
      port map(A => \temp_c6\, B => \temp[7]_net_1\, C => 
        \temp[8]_net_1\, Y => temp_n8);
    
    \pr_state_ns_a2_2[6]\ : NOR2A
      port map(A => CMOS_DrvX_0_SDramEn_0, B => 
        CMOS_DrvX_0_LVDSen_2, Y => \pr_state_ns_2[6]\);
    
    \temp[3]\ : DFN1E0C0
      port map(D => temp_n3, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => un2, Q => \temp[3]_net_1\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \pr_state_RNO_2[8]\ : OR3A
      port map(A => \pr_state[8]_net_1\, B => ref_ok_1, C => 
        ref_ok_2, Y => N_164);
    
    SD_RefEn_RNO : OR2
      port map(A => \pr_state[8]_net_1\, B => \pr_state[3]_net_1\, 
        Y => \SD_RefEn_RNO\);
    
    \pr_state_RNO[6]\ : AOI1B
      port map(A => N_160, B => N_159, C => \pr_state_ns_2[6]\, Y
         => \pr_state_ns[5]\);
    
    \pr_state_RNO[5]\ : NOR3C
      port map(A => \pr_state[11]_net_1\, B => SDram_rd_0_SD_RdOK, 
        C => \pr_state_ns_2[6]\, Y => \pr_state_ns[6]\);
    
    \pr_state[3]\ : DFN1C0
      port map(D => \pr_state_ns_i[8]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \pr_state[3]_net_1\);
    
    \temp[5]\ : DFN1E0C0
      port map(D => temp_n5, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => un2, Q => \temp[5]_net_1\);
    
    temp_n10_0 : XOR2
      port map(A => \temp_c9\, B => \temp[10]_net_1\, Y => 
        temp_n10);
    
    SD_wrEn_RNIVCK3 : INV
      port map(A => \Sdram_ctl_v2_0_SD_wrEn\, Y => 
        Sdram_ctl_v2_0_SD_wrEn_i);
    
    temp_c9 : NOR2A
      port map(A => \temp[9]_net_1\, B => \temp_c8\, Y => 
        \temp_c9\);
    
    \pr_state_RNO_1[9]\ : NOR2
      port map(A => \pr_state[9]_net_1\, B => Fifo_wr_0_AFULL, Y
         => N_175);
    
    \temp[1]\ : DFN1E0C0
      port map(D => temp_n1, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => un2, Q => \temp[1]_net_1\);
    
    SD_RefEn : DFN1C0
      port map(D => \SD_RefEn_RNO\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => Sdram_ctl_v2_0_SD_RefEn);
    
    temp_c8 : OR3B
      port map(A => \temp[7]_net_1\, B => \temp[8]_net_1\, C => 
        \temp_c6\, Y => \temp_c8\);
    
    \pr_state[2]\ : DFN1C0
      port map(D => \pr_state_RNO_0[2]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \pr_state[2]_net_1\);
    
    temp_n2_0 : AX1C
      port map(A => \temp[0]_net_1\, B => \temp[1]_net_1\, C => 
        \temp[2]_net_1\, Y => temp_n2);
    
    SD_rdEn_RNI2SH3 : INV
      port map(A => \Sdram_ctl_v2_0_SD_rdEn\, Y => 
        Sdram_ctl_v2_0_SD_rdEn_i);
    
    \pr_state_RNO[0]\ : NOR2B
      port map(A => \pr_state_ns[8]\, B => \pr_state[1]_net_1\, Y
         => \pr_state_RNO[0]_net_1\);
    
    \temp[2]\ : DFN1E0C0
      port map(D => temp_n2, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => un2, Q => \temp[2]_net_1\);
    
    \pr_state_ns_i_a2_0[0]\ : OR2
      port map(A => CMOS_DrvX_0_SDramEn_0, B => 
        CMOS_DrvX_0_LVDSen_2, Y => \pr_state_ns[8]\);
    
    \pr_state[7]\ : DFN1P0
      port map(D => \pr_state_RNO[7]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, PRE => PLL_Test1_0_SysRst_O, Q
         => \pr_state[7]_net_1\);
    
    \temp_RNIIRCF[2]\ : OA1
      port map(A => \temp[0]_net_1\, B => \temp[1]_net_1\, C => 
        \temp[2]_net_1\, Y => un2lt4);
    
    temp_10 : MX2
      port map(A => temp_n10, B => \temp[11]_net_1\, S => un2, Y
         => \temp_10\);
    
    temp_c2 : OR3C
      port map(A => \temp[0]_net_1\, B => \temp[1]_net_1\, C => 
        \temp[2]_net_1\, Y => \temp_c2\);
    
    PowerOK_RNO : OR2
      port map(A => un2, B => \SD_cke_c_c[0]\, Y => \PowerOK_RNO\);
    
    \pr_state_RNO_0[7]\ : NOR2A
      port map(A => \pr_state[7]_net_1\, B => 
        Sdram_ini_0_Sd_iniOK, Y => N_167);
    
    \temp_RNI4Q491[2]\ : OA1
      port map(A => un2lt4, B => un2lto4_0, C => un2lto7_1, Y => 
        un2lt9);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \pr_state_RNO_1[8]\ : AO1A
      port map(A => \pr_state_RNITULC[11]_net_1\, B => N_164, C
         => N_177, Y => \pr_state_ns_i_0[3]\);
    
    temp_c4 : OR3B
      port map(A => \temp[3]_net_1\, B => \temp[4]_net_1\, C => 
        \temp_c2\, Y => \temp_c4\);
    
    \pr_state_RNO[4]\ : NOR3A
      port map(A => \pr_state_ns[8]\, B => N_182, C => 
        \pr_state_ns_i_0[7]\, Y => \pr_state_RNO[4]_net_1\);
    
    \pr_state_RNO[1]\ : NOR2B
      port map(A => \pr_state_ns[8]\, B => \pr_state[2]_net_1\, Y
         => \pr_state_RNO_0[1]\);
    
    SD_rdEn : DFN1C0
      port map(D => \pr_state_RNITULC[11]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \Sdram_ctl_v2_0_SD_rdEn\);
    
    \pr_state_RNO[9]\ : NOR3A
      port map(A => \pr_state_ns[8]\, B => N_174, C => N_175, Y
         => \pr_state_RNO[9]_net_1\);
    
    \pr_state[0]\ : DFN1C0
      port map(D => \pr_state_RNO[0]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \pr_state[0]_net_1\);
    
    \pr_state_RNO[2]\ : NOR3B
      port map(A => \pr_state[4]_net_1\, B => \pr_state_ns[8]\, C
         => Fifo_rd_0_AFULL, Y => \pr_state_RNO_0[2]\);
    
    temp_20_0 : XNOR2
      port map(A => \temp[0]_net_1\, B => un2, Y => \temp_20_0\);
    
    \temp[6]\ : DFN1E0C0
      port map(D => temp_n6, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => un2, Q => \temp[6]_net_1\);
    
    \temp[11]\ : DFN1E0C0
      port map(D => temp_n11, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => un2, Q => \temp[11]_net_1\);
    
    \temp[8]\ : DFN1E0C0
      port map(D => temp_n8, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => un2, Q => \temp[8]_net_1\);
    
    \temp[0]\ : DFN1C0
      port map(D => \temp_20_0\, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \temp[0]_net_1\);
    
    PowerOK : DFN1C0
      port map(D => \PowerOK_RNO\, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \SD_cke_c_c[0]\);
    
    \temp_RNIH69A[4]\ : OR2
      port map(A => \temp[3]_net_1\, B => \temp[4]_net_1\, Y => 
        un2lto4_0);
    
    \temp[4]\ : DFN1E0C0
      port map(D => temp_n4, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => un2, Q => \temp[4]_net_1\);
    
    SD_pdEN : DFN1C0
      port map(D => \pr_state[3]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => Sdram_ctl_v2_0_SD_pdEN);
    
    \pr_state_RNO_0[8]\ : NOR3
      port map(A => \pr_state[8]_net_1\, B => 
        \pr_state[10]_net_1\, C => CMOS_DrvX_0_LVDSen_1, Y => 
        N_178);
    
    temp_n4_0 : AX1
      port map(A => \temp_c2\, B => \temp[3]_net_1\, C => 
        \temp[4]_net_1\, Y => temp_n4);
    
    \pr_state[9]\ : DFN1C0
      port map(D => \pr_state_RNO[9]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \pr_state[9]_net_1\);
    
    \pr_state[4]\ : DFN1C0
      port map(D => \pr_state_RNO[4]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \pr_state[4]_net_1\);
    
    \pr_state_RNO_4[4]\ : OR2
      port map(A => Sdram_ini_0_Sd_iniOK, B => 
        \pr_state[4]_net_1\, Y => \pr_state_ns_i_a2_0_0[7]\);
    
    \pr_state_RNO_2[4]\ : OR2
      port map(A => \pr_state[4]_net_1\, B => \pr_state[7]_net_1\, 
        Y => \pr_state_ns_i_a2_0[7]\);
    
    \temp_RNIREAA[8]\ : OR2
      port map(A => \temp[8]_net_1\, B => \temp[9]_net_1\, Y => 
        un2lto9_0);
    
    \pr_state_RNO_2[10]\ : NOR2B
      port map(A => \pr_state[9]_net_1\, B => SDRAM_wr_0_SD_WrOK, 
        Y => N_163);
    
    \pr_state_RNO[8]\ : NOR3A
      port map(A => \pr_state_ns[8]\, B => N_178, C => 
        \pr_state_ns_i_0[3]\, Y => \pr_state_RNO[8]_net_1\);
    
    \pr_state[6]\ : DFN1C0
      port map(D => \pr_state_ns[5]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \pr_state[6]_net_1\);
    
    \pr_state[10]\ : DFN1C0
      port map(D => \pr_state_RNO[10]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \pr_state[10]_net_1\);
    
    \pr_state_RNO_1[10]\ : NOR3A
      port map(A => SDram_rd_0_SD_RdOK, B => \pr_state[5]_net_1\, 
        C => \pr_state[9]_net_1\, Y => N_173);
    
    \pr_state_RNO_0[10]\ : NOR3
      port map(A => \pr_state[10]_net_1\, B => 
        \pr_state[5]_net_1\, C => N_163, Y => N_172);
    
    \pr_state_RNO[7]\ : OA1
      port map(A => N_167, B => \pr_state[3]_net_1\, C => 
        \pr_state_ns[8]\, Y => \pr_state_RNO[7]_net_1\);
    
    \pr_state_RNO[10]\ : NOR3A
      port map(A => \pr_state_ns[8]\, B => N_172, C => N_173, Y
         => \pr_state_RNO[10]_net_1\);
    
    temp_n7_0 : XNOR2
      port map(A => \temp_c6\, B => \temp[7]_net_1\, Y => temp_n7);
    
    \pr_state[8]\ : DFN1C0
      port map(D => \pr_state_RNO[8]_net_1\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \pr_state[8]_net_1\);
    
    \pr_state[1]\ : DFN1C0
      port map(D => \pr_state_RNO_0[1]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \pr_state[1]_net_1\);
    
    temp_n1_0 : XOR2
      port map(A => \temp[1]_net_1\, B => \temp[0]_net_1\, Y => 
        temp_n1);
    
    \pr_state_RNO_3[4]\ : OR2
      port map(A => \pr_state[7]_net_1\, B => Fifo_rd_0_AFULL, Y
         => \pr_state_ns_i_a2_1_0[7]\);
    
    \pr_state_RNITULC[11]\ : OR2
      port map(A => \pr_state[11]_net_1\, B => 
        \pr_state[10]_net_1\, Y => \pr_state_RNITULC[11]_net_1\);
    
    temp_n9_0 : XNOR2
      port map(A => \temp_c8\, B => \temp[9]_net_1\, Y => temp_n9);
    
    \pr_state_RNI1EA3[6]\ : OR2A
      port map(A => \pr_state[6]_net_1\, B => Fifo_wr_0_AFULL, Y
         => N_159);
    
    temp_n6_0 : AX1
      port map(A => \temp_c4\, B => \temp[5]_net_1\, C => 
        \temp[6]_net_1\, Y => temp_n6);
    
    \pr_state[5]\ : DFN1C0
      port map(D => \pr_state_ns[6]\, CLK => 
        PLL_Test1_0_Sys_66M_Clk, CLR => PLL_Test1_0_SysRst_O, Q
         => \pr_state[5]_net_1\);
    
    temp_n11_0 : AX1C
      port map(A => \temp[10]_net_1\, B => \temp_c9\, C => 
        \temp[11]_net_1\, Y => temp_n11);
    
    temp_c6 : OR3B
      port map(A => \temp[5]_net_1\, B => \temp[6]_net_1\, C => 
        \temp_c4\, Y => \temp_c6\);
    
    \pr_state_RNO_3[8]\ : NOR2
      port map(A => \pr_state[8]_net_1\, B => SDram_rd_0_SD_RdOK, 
        Y => N_177);
    
    \pr_state_RNO[3]\ : INV
      port map(A => \pr_state_ns[8]\, Y => \pr_state_ns_i[8]\);
    
    temp_n5_0 : XNOR2
      port map(A => \temp_c4\, B => \temp[5]_net_1\, Y => temp_n5);
    
    \pr_state_RNO_2[11]\ : NOR2A
      port map(A => CMOS_DrvX_0_LVDSen_2, B => N_159, Y => N_162);
    
    \temp[7]\ : DFN1E0C0
      port map(D => temp_n7, CLK => PLL_Test1_0_Sys_66M_Clk, CLR
         => PLL_Test1_0_SysRst_O, E => un2, Q => \temp[7]_net_1\);
    
    \pr_state_RNO_1[11]\ : NOR3A
      port map(A => SDram_rd_0_SD_RdOK, B => \pr_state[6]_net_1\, 
        C => \pr_state[0]_net_1\, Y => N_171);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    \temp[10]\ : DFN1C0
      port map(D => \temp_10\, CLK => PLL_Test1_0_Sys_66M_Clk, 
        CLR => PLL_Test1_0_SysRst_O, Q => \temp[10]_net_1\);
    
    \pr_state_RNO_0[11]\ : NOR3
      port map(A => \pr_state[11]_net_1\, B => 
        \pr_state[0]_net_1\, C => N_162, Y => N_169);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3;
use proasic3.all;

entity My_adder0_2 is

    port( intData2acc_RNI2KS7                         : in    std_logic_vector(28 to 28);
          intData2acc_RNI1KS7                         : in    std_logic_vector(27 to 27);
          intData2acc_RNI6JV9                         : in    std_logic_vector(33 to 33);
          intData2acc_RNI2BV9                         : in    std_logic_vector(18 to 18);
          intData2acc_RNI3BV9                         : in    std_logic_vector(19 to 19);
          intData2acc_RNIBN36                         : in    std_logic_vector(22 to 22);
          intData2acc_RNI3JV9                         : in    std_logic_vector(30 to 30);
          intData2acc_RNI5JV9                         : in    std_logic_vector(32 to 32);
          intData2acc_RNITEV9                         : in    std_logic_vector(20 to 20);
          intData2acc_RNIAN36                         : in    std_logic_vector(21 to 21);
          intData2acc_RNI4JV9                         : in    std_logic_vector(31 to 31);
          intData2acc_RNIDN36                         : in    std_logic_vector(24 to 24);
          intData2acc_RNIEN36                         : in    std_logic_vector(25 to 25);
          intData2acc_RNI9FV9                         : in    std_logic_vector(29 to 29);
          intData2acc_RNI8JV9                         : in    std_logic_vector(35 to 35);
          intData2acc_RNITJS7                         : in    std_logic_vector(23 to 23);
          intData2acc_RNI0KS7                         : in    std_logic_vector(26 to 26);
          intData2acc_RNI7JV9                         : in    std_logic_vector(34 to 34);
          \Z\\My_adder0_1_Sum_[15]\\\                 : out   std_logic;
          \Z\\My_adder0_1_Sum_[12]\\\                 : out   std_logic;
          \Z\\My_adder0_1_Sum_[6]\\\                  : out   std_logic;
          \Z\\My_adder0_1_Sum_[10]\\\                 : out   std_logic;
          \Z\\My_adder0_1_Sum_[9]\\\                  : out   std_logic;
          \Z\\My_adder0_1_Sum_[7]\\\                  : out   std_logic;
          \Z\\My_adder0_1_Sum_[11]\\\                 : out   std_logic;
          \Z\\My_adder0_1_Sum_[1]\\\                  : out   std_logic;
          \Z\\My_adder0_1_Sum_[3]\\\                  : out   std_logic;
          \Z\\My_adder0_1_Sum_[13]\\\                 : out   std_logic;
          \Z\\adc_muxtmp_test_0_DataOut27to14_[14]\\\ : in    std_logic;
          \Z\\My_adder0_1_Sum_[0]\\\                  : out   std_logic;
          \Z\\My_adder0_1_Sum_[8]\\\                  : out   std_logic;
          \Z\\My_adder0_1_Sum_[14]\\\                 : out   std_logic;
          \Z\\My_adder0_1_Sum_[2]\\\                  : out   std_logic;
          \Z\\My_adder0_1_Sum_[4]\\\                  : out   std_logic;
          \Z\\My_adder0_1_Sum_[5]\\\                  : out   std_logic;
          \Z\\My_adder0_1_Sum_[17]\\\                 : out   std_logic;
          My_adder0_2_GND                             : in    std_logic;
          \Z\\My_adder0_1_Sum_[16]\\\                 : out   std_logic
        );

end My_adder0_2;

architecture DEF_ARCH of My_adder0_2 is 

  component XOR3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component MAJ3
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          C : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component AND2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

  component XOR2
    port( A : in    std_logic := 'U';
          B : in    std_logic := 'U';
          Y : out   std_logic
        );
  end component;

    signal Carry_15_net, Carry_8_net, Carry_7_net, Carry_5_net, 
        Carry_4_net, Carry_16_net, Carry_11_net, Carry_10_net, 
        Carry_6_net, Carry_13_net, Carry_12_net, Carry_3_net, 
        Carry_2_net, Carry_1_net, Carry_14_net, Carry_0_net, 
        Carry_9_net, \GND\, \VCC\, GND_0, VCC_0 : std_logic;

begin 


    XOR3_Sum_16_inst : XOR3
      port map(A => My_adder0_2_GND, B => intData2acc_RNI7JV9(34), 
        C => Carry_15_net, Y => \Z\\My_adder0_1_Sum_[16]\\\);
    
    MAJ3_Carry_8_inst : MAJ3
      port map(A => Carry_7_net, B => My_adder0_2_GND, C => 
        intData2acc_RNI0KS7(26), Y => Carry_8_net);
    
    MAJ3_Carry_9_inst : MAJ3
      port map(A => Carry_8_net, B => My_adder0_2_GND, C => 
        intData2acc_RNI1KS7(27), Y => Carry_9_net);
    
    XOR3_Sum_5_inst : XOR3
      port map(A => My_adder0_2_GND, B => intData2acc_RNITJS7(23), 
        C => Carry_4_net, Y => \Z\\My_adder0_1_Sum_[5]\\\);
    
    XOR3_Sum_2_inst : XOR3
      port map(A => My_adder0_2_GND, B => intData2acc_RNITEV9(20), 
        C => Carry_1_net, Y => \Z\\My_adder0_1_Sum_[2]\\\);
    
    XOR3_Sum_4_inst : XOR3
      port map(A => My_adder0_2_GND, B => intData2acc_RNIBN36(22), 
        C => Carry_3_net, Y => \Z\\My_adder0_1_Sum_[4]\\\);
    
    XOR3_Sum_11_inst : XOR3
      port map(A => My_adder0_2_GND, B => intData2acc_RNI9FV9(29), 
        C => Carry_10_net, Y => \Z\\My_adder0_1_Sum_[11]\\\);
    
    XOR3_Sum_12_inst : XOR3
      port map(A => My_adder0_2_GND, B => intData2acc_RNI3JV9(30), 
        C => Carry_11_net, Y => \Z\\My_adder0_1_Sum_[12]\\\);
    
    MAJ3_Carry_5_inst : MAJ3
      port map(A => Carry_4_net, B => My_adder0_2_GND, C => 
        intData2acc_RNITJS7(23), Y => Carry_5_net);
    
    MAJ3_Carry_2_inst : MAJ3
      port map(A => Carry_1_net, B => My_adder0_2_GND, C => 
        intData2acc_RNITEV9(20), Y => Carry_2_net);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    MAJ3_Carry_1_inst : MAJ3
      port map(A => Carry_0_net, B => My_adder0_2_GND, C => 
        intData2acc_RNI3BV9(19), Y => Carry_1_net);
    
    MAJ3_Carry_4_inst : MAJ3
      port map(A => Carry_3_net, B => My_adder0_2_GND, C => 
        intData2acc_RNIBN36(22), Y => Carry_4_net);
    
    XOR3_Sum_13_inst : XOR3
      port map(A => My_adder0_2_GND, B => intData2acc_RNI4JV9(31), 
        C => Carry_12_net, Y => \Z\\My_adder0_1_Sum_[13]\\\);
    
    XOR3_Sum_1_inst : XOR3
      port map(A => My_adder0_2_GND, B => intData2acc_RNI3BV9(19), 
        C => Carry_0_net, Y => \Z\\My_adder0_1_Sum_[1]\\\);
    
    MAJ3_Carry_12_inst : MAJ3
      port map(A => Carry_11_net, B => My_adder0_2_GND, C => 
        intData2acc_RNI3JV9(30), Y => Carry_12_net);
    
    XOR3_Sum_17_inst : XOR3
      port map(A => My_adder0_2_GND, B => intData2acc_RNI8JV9(35), 
        C => Carry_16_net, Y => \Z\\My_adder0_1_Sum_[17]\\\);
    
    MAJ3_Carry_7_inst : MAJ3
      port map(A => Carry_6_net, B => My_adder0_2_GND, C => 
        intData2acc_RNIEN36(25), Y => Carry_7_net);
    
    GND_i : GND
      port map(Y => \GND\);
    
    XOR3_Sum_6_inst : XOR3
      port map(A => My_adder0_2_GND, B => intData2acc_RNIDN36(24), 
        C => Carry_5_net, Y => \Z\\My_adder0_1_Sum_[6]\\\);
    
    MAJ3_Carry_14_inst : MAJ3
      port map(A => Carry_13_net, B => My_adder0_2_GND, C => 
        intData2acc_RNI5JV9(32), Y => Carry_14_net);
    
    MAJ3_Carry_13_inst : MAJ3
      port map(A => Carry_12_net, B => My_adder0_2_GND, C => 
        intData2acc_RNI4JV9(31), Y => Carry_13_net);
    
    XOR3_Sum_3_inst : XOR3
      port map(A => My_adder0_2_GND, B => intData2acc_RNIAN36(21), 
        C => Carry_2_net, Y => \Z\\My_adder0_1_Sum_[3]\\\);
    
    XOR3_Sum_14_inst : XOR3
      port map(A => My_adder0_2_GND, B => intData2acc_RNI5JV9(32), 
        C => Carry_13_net, Y => \Z\\My_adder0_1_Sum_[14]\\\);
    
    XOR3_Sum_8_inst : XOR3
      port map(A => My_adder0_2_GND, B => intData2acc_RNI0KS7(26), 
        C => Carry_7_net, Y => \Z\\My_adder0_1_Sum_[8]\\\);
    
    MAJ3_Carry_11_inst : MAJ3
      port map(A => Carry_10_net, B => My_adder0_2_GND, C => 
        intData2acc_RNI9FV9(29), Y => Carry_11_net);
    
    MAJ3_Carry_16_inst : MAJ3
      port map(A => Carry_15_net, B => My_adder0_2_GND, C => 
        intData2acc_RNI7JV9(34), Y => Carry_16_net);
    
    XOR3_Sum_7_inst : XOR3
      port map(A => My_adder0_2_GND, B => intData2acc_RNIEN36(25), 
        C => Carry_6_net, Y => \Z\\My_adder0_1_Sum_[7]\\\);
    
    MAJ3_Carry_10_inst : MAJ3
      port map(A => Carry_9_net, B => My_adder0_2_GND, C => 
        intData2acc_RNI2KS7(28), Y => Carry_10_net);
    
    MAJ3_Carry_3_inst : MAJ3
      port map(A => Carry_2_net, B => My_adder0_2_GND, C => 
        intData2acc_RNIAN36(21), Y => Carry_3_net);
    
    XOR3_Sum_15_inst : XOR3
      port map(A => My_adder0_2_GND, B => intData2acc_RNI6JV9(33), 
        C => Carry_14_net, Y => \Z\\My_adder0_1_Sum_[15]\\\);
    
    AND2_Carry_0_inst : AND2
      port map(A => \Z\\adc_muxtmp_test_0_DataOut27to14_[14]\\\, 
        B => intData2acc_RNI2BV9(18), Y => Carry_0_net);
    
    MAJ3_Carry_15_inst : MAJ3
      port map(A => Carry_14_net, B => My_adder0_2_GND, C => 
        intData2acc_RNI6JV9(33), Y => Carry_15_net);
    
    XOR3_Sum_9_inst : XOR3
      port map(A => My_adder0_2_GND, B => intData2acc_RNI1KS7(27), 
        C => Carry_8_net, Y => \Z\\My_adder0_1_Sum_[9]\\\);
    
    XOR2_Sum_0_inst : XOR2
      port map(A => \Z\\adc_muxtmp_test_0_DataOut27to14_[14]\\\, 
        B => intData2acc_RNI2BV9(18), Y => 
        \Z\\My_adder0_1_Sum_[0]\\\);
    
    MAJ3_Carry_6_inst : MAJ3
      port map(A => Carry_5_net, B => My_adder0_2_GND, C => 
        intData2acc_RNIDN36(24), Y => Carry_6_net);
    
    XOR3_Sum_10_inst : XOR3
      port map(A => My_adder0_2_GND, B => intData2acc_RNI2KS7(28), 
        C => Carry_9_net, Y => \Z\\My_adder0_1_Sum_[10]\\\);
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    

end DEF_ARCH; 

library ieee;
use ieee.std_logic_1164.all;
library proasic3;
use proasic3.all;

entity smart_top is

    port( ExterCLk    : in    std_logic;
          CMOS_sample : out   std_logic;
          mem_HL      : out   std_logic;
          Sync_X      : out   std_logic;
          Clock_Y     : out   std_logic;
          spi_data    : out   std_logic;
          reset_ds    : out   std_logic;
          Clock_X     : out   std_logic;
          Prebus1     : out   std_logic;
          Prebus2     : out   std_logic;
          Sync_Y      : out   std_logic;
          spi_clock   : out   std_logic;
          Sh_co       : out   std_logic;
          precharge   : out   std_logic;
          AdcClk      : out   std_logic;
          VoltAvg     : out   std_logic;
          NoRowSel    : out   std_logic;
          CMOS_reset  : out   std_logic;
          Pre_co      : out   std_logic;
          spi_load    : out   std_logic;
          SD_ras_n    : out   std_logic;
          SD_cas_n    : out   std_logic;
          SD_we_n     : out   std_logic;
          LVDS_O      : out   std_logic;
          tok         : out   std_logic;
          DRY         : out   std_logic;
          Sd_DQ       : inout std_logic_vector(71 downto 0) := (others => 'Z');
          SD_cke      : out   std_logic_vector(1 downto 0);
          SD_cs_n     : out   std_logic_vector(1 downto 0);
          SD_Clk      : out   std_logic_vector(1 downto 0);
          SD_dqm      : out   std_logic_vector(7 downto 0);
          SD_addr     : out   std_logic_vector(12 downto 0);
          SD_ba       : out   std_logic_vector(1 downto 0);
          ADCdataIn   : in    std_logic_vector(13 downto 0)
        );

end smart_top;

architecture DEF_ARCH of smart_top is 

  component BIBUF
    port( PAD : inout   std_logic;
          D   : in    std_logic := 'U';
          E   : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component OUTBUF
    port( D   : in    std_logic := 'U';
          PAD : out   std_logic
        );
  end component;

  component FrameMk
    port( FrameMk_GND             : in    std_logic := 'U';
          CMOS_DrvX_0_LVDSen_3    : in    std_logic := 'U';
          FrameMk_VCC             : in    std_logic := 'U';
          CMOS_DrvX_0_LVDSen      : in    std_logic := 'U';
          tok_c                   : out   std_logic;
          LVDS_O_c                : out   std_logic;
          Main_ctl4SD_0_ByteRdEn  : in    std_logic := 'U';
          CMOS_DrvX_0_LVDSen_2    : in    std_logic := 'U';
          CMOS_DrvX_0_LVDSen_1    : in    std_logic := 'U';
          CMOS_DrvX_0_LVDSen_0    : in    std_logic := 'U';
          FrameMk_0_LVDS_ok       : out   std_logic;
          FrameMk_0_LVDS_ok_i     : out   std_logic;
          PLL_Test1_0_SysRst_O    : in    std_logic := 'U';
          PLL_Test1_0_Sys_66M_Clk : in    std_logic := 'U'
        );
  end component;

  component My_adder0_1
    port( intData2acc_RNIEVV9                         : in    std_logic_vector(64 to 64) := (others => 'U');
          intData2acc_RNIDVV9                         : in    std_logic_vector(63 to 63) := (others => 'U');
          intData2acc_RNIGVV9                         : in    std_logic_vector(66 to 66) := (others => 'U');
          intData2acc_RNIDRV9                         : in    std_logic_vector(56 to 56) := (others => 'U');
          intData2acc_RNIERV9                         : in    std_logic_vector(57 to 57) := (others => 'U');
          intData2acc_RNIHVV9                         : in    std_logic_vector(67 to 67) := (others => 'U');
          intData2acc_RNIAVV9                         : in    std_logic_vector(60 to 60) := (others => 'U');
          intData2acc_RNIBVV9                         : in    std_logic_vector(61 to 61) := (others => 'U');
          intData2acc_RNIFVV9                         : in    std_logic_vector(65 to 65) := (others => 'U');
          intData2acc_RNIPB46                         : in    std_logic_vector(71 to 71) := (others => 'U');
          intData2acc_RNIGRV9                         : in    std_logic_vector(59 downto 58) := (others => 'U');
          intData2acc_RNICVV9                         : in    std_logic_vector(62 to 62) := (others => 'U');
          intData2acc_RNID30A                         : in    std_logic_vector(70 to 70) := (others => 'U');
          intData2acc_RNIARV9                         : in    std_logic_vector(54 to 54) := (others => 'U');
          intData2acc_RNIBRV9                         : in    std_logic_vector(55 to 55) := (others => 'U');
          \Z\\My_adder0_3_Sum_[15]\\\                 : out   std_logic;
          \Z\\My_adder0_3_Sum_[12]\\\                 : out   std_logic;
          \Z\\My_adder0_3_Sum_[6]\\\                  : out   std_logic;
          \Z\\My_adder0_3_Sum_[10]\\\                 : out   std_logic;
          \Z\\My_adder0_3_Sum_[9]\\\                  : out   std_logic;
          \Z\\My_adder0_3_Sum_[7]\\\                  : out   std_logic;
          N_6                                         : in    std_logic := 'U';
          \Z\\My_adder0_3_Sum_[11]\\\                 : out   std_logic;
          \Z\\My_adder0_3_Sum_[1]\\\                  : out   std_logic;
          \Z\\My_adder0_3_Sum_[3]\\\                  : out   std_logic;
          \Z\\My_adder0_3_Sum_[13]\\\                 : out   std_logic;
          \Z\\My_adder0_3_Sum_[0]\\\                  : out   std_logic;
          \Z\\My_adder0_3_Sum_[8]\\\                  : out   std_logic;
          \Z\\My_adder0_3_Sum_[14]\\\                 : out   std_logic;
          \Z\\My_adder0_3_Sum_[2]\\\                  : out   std_logic;
          \Z\\My_adder0_3_Sum_[4]\\\                  : out   std_logic;
          N_4                                         : in    std_logic := 'U';
          \Z\\My_adder0_3_Sum_[5]\\\                  : out   std_logic;
          \Z\\My_adder0_3_Sum_[17]\\\                 : out   std_logic;
          My_adder0_1_GND                             : in    std_logic := 'U';
          \Z\\My_adder0_3_Sum_[16]\\\                 : out   std_logic;
          \Z\\adc_muxtmp_test_0_DataOut55to42_[43]\\\ : in    std_logic := 'U'
        );
  end component;

  component Fifo_rd
    port( \Z\\Fifo_wr_0_Q_[27]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[23]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[69]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[1]\\\              : out   std_logic;
          \Z\\Fifo_wr_0_Q_[67]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[4]\\\              : out   std_logic;
          \Z\\Fifo_wr_0_Q_[63]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[7]\\\              : out   std_logic;
          \Z\\Fifo_wr_0_Q_[56]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[25]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[24]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[48]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[65]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[64]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[51]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[38]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[71]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[50]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[70]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[18]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[6]\\\              : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[71]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[70]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[69]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[68]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[67]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[66]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[65]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[64]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[63]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[62]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[61]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[60]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[59]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[58]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[57]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[56]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[55]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[54]\\\ : in    std_logic := 'U';
          \Z\\Fifo_wr_0_Q_[46]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[52]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[36]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[59]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[0]\\\              : out   std_logic;
          \Z\\Fifo_wr_0_Q_[16]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[57]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[41]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[53]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[40]\\\             : out   std_logic;
          Sdram_cmd_0_WFifo_re                : in    std_logic := 'U';
          \Z\\Fifo_wr_0_Q_[31]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[28]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[30]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[42]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[11]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[10]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[55]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[68]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[54]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[49]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[9]\\\              : out   std_logic;
          \Z\\Fifo_wr_0_Q_[5]\\\              : out   std_logic;
          Fifo_wr_0_AFULL                     : out   std_logic;
          \Z\\Fifo_wr_0_Q_[32]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[47]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[43]\\\             : out   std_logic;
          Main_ctl4SD_0_fifo_rst_n_3          : in    std_logic := 'U';
          \Z\\Fifo_wr_0_Q_[12]\\\             : out   std_logic;
          Main_ctl4SD_0_Fifo_wr               : in    std_logic := 'U';
          \Z\\Fifo_wr_0_Q_[26]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[39]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[19]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[37]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[3]\\\              : out   std_logic;
          \Z\\Fifo_wr_0_Q_[33]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[66]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[17]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[13]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[45]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[44]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[21]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[2]\\\              : out   std_logic;
          \Z\\Fifo_wr_0_Q_[20]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[61]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[35]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[34]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[60]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[15]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[14]\\\             : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[35]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[34]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[33]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[32]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[31]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[30]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[29]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[28]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[27]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[26]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[25]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[24]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[23]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[22]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[21]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[20]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[19]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[18]\\\ : in    std_logic := 'U';
          Main_ctl4SD_0_fifo_rst_n_4          : in    std_logic := 'U';
          \Z\\Fifo_wr_0_Q_[22]\\\             : out   std_logic;
          \Z\\Fifo_wr_0_Q_[8]\\\              : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[53]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[52]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[51]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[50]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[49]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[48]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[47]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[46]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[45]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[44]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[43]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[42]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[41]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[40]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[39]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[38]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[37]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[36]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[17]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[16]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[15]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[14]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[13]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[12]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[11]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[10]\\\ : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[9]\\\  : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[8]\\\  : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[7]\\\  : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[6]\\\  : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[5]\\\  : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[4]\\\  : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[3]\\\  : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[2]\\\  : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[1]\\\  : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[0]\\\  : in    std_logic := 'U';
          Fifo_rd_VCC                         : in    std_logic := 'U';
          Main_ctl4SD_0_fifo_rst_n            : in    std_logic := 'U';
          \Z\\Fifo_wr_0_Q_[62]\\\             : out   std_logic;
          Main_ctl4SD_0_fifo_rst_n_5          : in    std_logic := 'U';
          \Z\\Fifo_wr_0_Q_[29]\\\             : out   std_logic;
          Main_ctl4SD_0_fifo_rst_n_6          : in    std_logic := 'U';
          PLL_Test1_0_Sys_66M_Clk             : in    std_logic := 'U';
          \Z\\Fifo_wr_0_Q_[58]\\\             : out   std_logic;
          Fifo_rd_GND                         : in    std_logic := 'U'
        );
  end component;

  component CMOS_DrvX
    port( CMOS_reset_c             : out   std_logic;
          CMOS_sample_c            : out   std_logic;
          precharge_c              : out   std_logic;
          mem_HL_c                 : out   std_logic;
          spi_load_c               : out   std_logic;
          spi_data_c               : out   std_logic;
          spi_clock_c              : out   std_logic;
          CMOS_DrvX_VCC            : in    std_logic := 'U';
          PLL_Test1_0_ADC_66M_Clk  : in    std_logic := 'U';
          DRY_c_c                  : out   std_logic;
          CMOS_DrvX_0_AdcEn        : out   std_logic;
          Sync_Y_c                 : out   std_logic;
          Clock_Y_c                : out   std_logic;
          NoRowSel_c               : out   std_logic;
          Pre_co_c                 : out   std_logic;
          Sh_co_c                  : out   std_logic;
          Sync_X_c                 : out   std_logic;
          Clock_X_c                : out   std_logic;
          CMOS_DrvX_0_LVDSen_3     : out   std_logic;
          PLL_Test1_0_Sys_66M_Clk  : in    std_logic := 'U';
          PLL_Test1_0_SysRst_O     : in    std_logic := 'U';
          CMOS_DrvX_0_LVDSen_2     : out   std_logic;
          CMOS_DrvX_0_LVDSen_1     : out   std_logic;
          CMOS_DrvX_0_LVDSen_0     : out   std_logic;
          CMOS_DrvX_0_SDramEn_5    : out   std_logic;
          CMOS_DrvX_0_SDramEn_4    : out   std_logic;
          CMOS_DrvX_0_SDramEn_3    : out   std_logic;
          CMOS_DrvX_0_SDramEn_2    : out   std_logic;
          CMOS_DrvX_0_SDramEn_1    : out   std_logic;
          CMOS_DrvX_0_SDramEn_0    : out   std_logic;
          Sdram_cmd_0_SDoneFrameOk : in    std_logic := 'U';
          FrameMk_0_LVDS_ok        : in    std_logic := 'U';
          CMOS_DrvX_0_LVDSen       : out   std_logic;
          CMOS_DrvX_0_SDramEn      : out   std_logic;
          CMOS_DrvX_GND            : in    std_logic := 'U'
        );
  end component;

  component My_adder0
    port( intData2acc_RNICNV9                         : in    std_logic_vector(46 to 46) := (others => 'U');
          intData2acc_RNIBNV9                         : in    std_logic_vector(45 to 45) := (others => 'U');
          intData2acc_RNI9RV9                         : in    std_logic_vector(51 to 51) := (others => 'U');
          intData2acc_RNI6JV9                         : in    std_logic_vector(36 to 36) := (others => 'U');
          intData2acc_RNI7JV9                         : in    std_logic_vector(37 to 37) := (others => 'U');
          intData2acc_RNI6NV9                         : in    std_logic_vector(40 to 40) := (others => 'U');
          intData2acc_RNIENV9                         : in    std_logic_vector(48 to 48) := (others => 'U');
          intData2acc_RNI8RV9                         : in    std_logic_vector(50 to 50) := (others => 'U');
          intData2acc_RNIBJV9                         : in    std_logic_vector(38 to 38) := (others => 'U');
          intData2acc_RNICJV9                         : in    std_logic_vector(39 to 39) := (others => 'U');
          intData2acc_RNIFNV9                         : in    std_logic_vector(49 to 49) := (others => 'U');
          intData2acc_RNI8NV9                         : in    std_logic_vector(42 to 42) := (others => 'U');
          intData2acc_RNI9NV9                         : in    std_logic_vector(43 to 43) := (others => 'U');
          intData2acc_RNIDNV9                         : in    std_logic_vector(47 to 47) := (others => 'U');
          intData2acc_RNI7NV9                         : in    std_logic_vector(41 to 41) := (others => 'U');
          intData2acc_RNIANV9                         : in    std_logic_vector(44 to 44) := (others => 'U');
          intData2acc_RNIBRV9                         : in    std_logic_vector(53 downto 52) := (others => 'U');
          \Z\\My_adder0_2_Sum_[15]\\\                 : out   std_logic;
          \Z\\My_adder0_2_Sum_[12]\\\                 : out   std_logic;
          \Z\\My_adder0_2_Sum_[6]\\\                  : out   std_logic;
          \Z\\My_adder0_2_Sum_[10]\\\                 : out   std_logic;
          \Z\\My_adder0_2_Sum_[9]\\\                  : out   std_logic;
          \Z\\My_adder0_2_Sum_[7]\\\                  : out   std_logic;
          \Z\\My_adder0_2_Sum_[11]\\\                 : out   std_logic;
          \Z\\My_adder0_2_Sum_[1]\\\                  : out   std_logic;
          \Z\\My_adder0_2_Sum_[3]\\\                  : out   std_logic;
          \Z\\My_adder0_2_Sum_[13]\\\                 : out   std_logic;
          \Z\\My_adder0_2_Sum_[0]\\\                  : out   std_logic;
          \Z\\My_adder0_2_Sum_[8]\\\                  : out   std_logic;
          \Z\\My_adder0_2_Sum_[14]\\\                 : out   std_logic;
          \Z\\adc_muxtmp_test_0_DataOut41to28_[29]\\\ : in    std_logic := 'U';
          \Z\\My_adder0_2_Sum_[2]\\\                  : out   std_logic;
          \Z\\My_adder0_2_Sum_[4]\\\                  : out   std_logic;
          \Z\\My_adder0_2_Sum_[5]\\\                  : out   std_logic;
          \Z\\My_adder0_2_Sum_[17]\\\                 : out   std_logic;
          My_adder0_GND                               : in    std_logic := 'U';
          \Z\\My_adder0_2_Sum_[16]\\\                 : out   std_logic
        );
  end component;

  component GND
    port( Y : out   std_logic
        );
  end component;

  component VCC
    port( Y : out   std_logic
        );
  end component;

  component INBUF
    port( PAD : in    std_logic := 'U';
          Y   : out   std_logic
        );
  end component;

  component SDRAM_wr
    port( \Z\\SDRAM_wr_0_wr_state_[2]\\\ : out   std_logic;
          \Z\\SDRAM_wr_0_wr_state_[1]\\\ : out   std_logic;
          \Z\\SDRAM_wr_0_wr_state_[0]\\\ : out   std_logic;
          Sdram_ctl_v2_0_SD_wrEn_i       : in    std_logic := 'U';
          PLL_Test1_0_SysRst_O           : in    std_logic := 'U';
          PLL_Test1_0_Sys_66M_Clk        : in    std_logic := 'U';
          SDRAM_wr_0_SD_WrOK             : out   std_logic;
          Sdram_cmd_0_wrrow_end          : in    std_logic := 'U';
          Sdram_ctl_v2_0_SD_wrEn         : in    std_logic := 'U'
        );
  end component;

  component Counter_ref
    port( refenlto5               : out   std_logic;
          Sdram_ctl_v2_0_SD_RefEn : in    std_logic := 'U';
          PLL_Test1_0_SysRst_O    : in    std_logic := 'U';
          PLL_Test1_0_Sys_66M_Clk : in    std_logic := 'U';
          Main_ctl4SD_0_ByteRdEn  : in    std_logic := 'U';
          CMOS_DrvX_0_LVDSen_2    : in    std_logic := 'U'
        );
  end component;

  component My_adder0_3
    port( intData2acc_RNI6J36         : in    std_logic_vector(10 to 10) := (others => 'U');
          intData2acc_RNIK507         : in    std_logic_vector(9 to 9) := (others => 'U');
          intData2acc_RNIBJ36         : in    std_logic_vector(15 to 15) := (others => 'U');
          intData2acc_RNIVOQA         : in    std_logic_vector(0 to 0) := (others => 'U');
          intData2acc_RNI0TQA         : in    std_logic_vector(1 to 1) := (others => 'U');
          intData2acc_RNIFHV6         : in    std_logic_vector(4 to 4) := (others => 'U');
          intData2acc_RNI8J36         : in    std_logic_vector(12 to 12) := (others => 'U');
          intData2acc_RNIAJ36         : in    std_logic_vector(14 to 14) := (others => 'U');
          intData2acc_RNI11RA         : in    std_logic_vector(2 to 2) := (others => 'U');
          intData2acc_RNIEDV6         : in    std_logic_vector(3 to 3) := (others => 'U');
          intData2acc_RNI9J36         : in    std_logic_vector(13 to 13) := (others => 'U');
          intData2acc_RNIHPV6         : in    std_logic_vector(6 to 6) := (others => 'U');
          intData2acc_RNIITV6         : in    std_logic_vector(7 to 7) := (others => 'U');
          intData2acc_RNI7J36         : in    std_logic_vector(11 to 11) := (others => 'U');
          intData2acc_RNIDJ36         : in    std_logic_vector(17 to 17) := (others => 'U');
          intData2acc_RNIGLV6         : in    std_logic_vector(5 to 5) := (others => 'U');
          intData2acc_RNIJ107         : in    std_logic_vector(8 to 8) := (others => 'U');
          intData2acc_RNICJ36         : in    std_logic_vector(16 to 16) := (others => 'U');
          \Z\\My_adder0_0_Sum_[15]\\\ : out   std_logic;
          \Z\\My_adder0_0_Sum_[12]\\\ : out   std_logic;
          \Z\\My_adder0_0_Sum_[6]\\\  : out   std_logic;
          \Z\\My_adder0_0_Sum_[10]\\\ : out   std_logic;
          \Z\\My_adder0_0_Sum_[9]\\\  : out   std_logic;
          \Z\\My_adder0_0_Sum_[7]\\\  : out   std_logic;
          \Z\\My_adder0_0_Sum_[11]\\\ : out   std_logic;
          \Z\\My_adder0_0_Sum_[1]\\\  : out   std_logic;
          \Z\\My_adder0_0_Sum_[3]\\\  : out   std_logic;
          \Z\\My_adder0_0_Sum_[13]\\\ : out   std_logic;
          \Z\\My_adder0_0_Sum_[0]\\\  : out   std_logic;
          \Z\\My_adder0_0_Sum_[8]\\\  : out   std_logic;
          \Z\\My_adder0_0_Sum_[14]\\\ : out   std_logic;
          \Z\\My_adder0_0_Sum_[2]\\\  : out   std_logic;
          \Z\\My_adder0_0_Sum_[4]\\\  : out   std_logic;
          \Z\\My_adder0_0_Sum_[5]\\\  : out   std_logic;
          \Z\\My_adder0_0_Sum_[17]\\\ : out   std_logic;
          My_adder0_3_GND             : in    std_logic := 'U';
          \Z\\My_adder0_0_Sum_[16]\\\ : out   std_logic
        );
  end component;

  component SDRAM_Ref
    port( \Z\\SDRAM_Ref_0_Ref_state_[2]\\\ : out   std_logic;
          \Z\\SDRAM_Ref_0_Ref_state_[1]\\\ : out   std_logic;
          \Z\\SDRAM_Ref_0_Ref_state_[0]\\\ : out   std_logic;
          ref_ok_1                         : out   std_logic;
          PLL_Test1_0_SysRst_O             : in    std_logic := 'U';
          PLL_Test1_0_Sys_66M_Clk          : in    std_logic := 'U';
          ref_ok_2                         : out   std_logic;
          Sdram_ctl_v2_0_SD_RefEn          : in    std_logic := 'U';
          Sdram_ini_0_Sd_iniOK             : in    std_logic := 'U';
          refenlto5                        : in    std_logic := 'U';
          Sdram_ctl_v2_0_SD_pdEN           : in    std_logic := 'U'
        );
  end component;

  component Sdram_cmd
    port( SD_cs_n_c_c                      : out   std_logic_vector(1 to 1);
          SD_dqm_c_c_c_c_c_c_c_c           : out   std_logic_vector(1 to 1);
          SD_cke_c_c                       : in    std_logic_vector(0 to 0) := (others => 'U');
          SD_Clk_c_c                       : out   std_logic_vector(1 to 1);
          SD_addr_c                        : out   std_logic_vector(12 downto 0);
          Sdram_cmd_0_RFifo_we             : out   std_logic;
          Sdram_cmd_0_rdrow_end            : out   std_logic;
          Sdram_cmd_0_WFifo_re             : out   std_logic;
          Sdram_cmd_0_wrrow_end            : out   std_logic;
          SD_ras_n_c                       : out   std_logic;
          SD_we_n_c                        : out   std_logic;
          SD_cas_n_c                       : out   std_logic;
          CMOS_DrvX_0_LVDSen               : in    std_logic := 'U';
          Sdram_cmd_0_SDoneFrameOk         : out   std_logic;
          CMOS_DrvX_0_SDramEn              : in    std_logic := 'U';
          PLL_Test1_0_SysRst_O             : in    std_logic := 'U';
          PLL_Test1_0_Sys_66M_Clk          : in    std_logic := 'U';
          LVDS_enReg                       : out   std_logic;
          CMOS_DrvX_0_LVDSen_2             : in    std_logic := 'U';
          \Z\\Sdram_ini_0_ini_state_[0]\\\ : in    std_logic := 'U';
          un6_sdramenreg                   : in    std_logic := 'U';
          N_264                            : out   std_logic;
          \Z\\SDRAM_Ref_0_Ref_state_[0]\\\ : in    std_logic := 'U';
          \Z\\SDRAM_Ref_0_Ref_state_[2]\\\ : in    std_logic := 'U';
          \Z\\SDRAM_Ref_0_Ref_state_[1]\\\ : in    std_logic := 'U';
          PLL_Test1_0_Sdram_clk            : in    std_logic := 'U';
          \Z\\SDram_rd_0_rd_state_[1]\\\   : in    std_logic := 'U';
          \Z\\SDram_rd_0_rd_state_[2]\\\   : in    std_logic := 'U';
          \Z\\SDram_rd_0_rd_state_[0]\\\   : in    std_logic := 'U';
          \Z\\Sdram_ini_0_ini_state_[2]\\\ : in    std_logic := 'U';
          \Z\\Sdram_ini_0_ini_state_[1]\\\ : in    std_logic := 'U';
          N_264_0                          : out   std_logic;
          N_264_1                          : out   std_logic;
          \Z\\SDRAM_wr_0_wr_state_[1]\\\   : in    std_logic := 'U';
          \Z\\SDRAM_wr_0_wr_state_[0]\\\   : in    std_logic := 'U';
          \Z\\SDRAM_wr_0_wr_state_[2]\\\   : in    std_logic := 'U';
          N_264_2                          : out   std_logic
        );
  end component;

  component Sdram_ini
    port( \Z\\Sdram_ini_0_ini_state_[2]\\\ : out   std_logic;
          \Z\\Sdram_ini_0_ini_state_[1]\\\ : out   std_logic;
          \Z\\Sdram_ini_0_ini_state_[0]\\\ : out   std_logic;
          PLL_Test1_0_SysRst_O             : in    std_logic := 'U';
          PLL_Test1_0_Sys_66M_Clk          : in    std_logic := 'U';
          Sdram_ctl_v2_0_SD_iniEn          : in    std_logic := 'U';
          Sdram_ini_0_Sd_iniOK             : out   std_logic;
          Sdram_ini_0_Sd_iniOK_i           : out   std_logic
        );
  end component;

  component SDram_rd
    port( \Z\\SDram_rd_0_rd_state_[2]\\\ : out   std_logic;
          \Z\\SDram_rd_0_rd_state_[1]\\\ : out   std_logic;
          \Z\\SDram_rd_0_rd_state_[0]\\\ : out   std_logic;
          Sdram_ctl_v2_0_SD_rdEn_i       : in    std_logic := 'U';
          PLL_Test1_0_SysRst_O           : in    std_logic := 'U';
          PLL_Test1_0_Sys_66M_Clk        : in    std_logic := 'U';
          SDram_rd_0_SD_RdOK             : out   std_logic;
          Sdram_ctl_v2_0_SD_rdEn         : in    std_logic := 'U';
          Sdram_cmd_0_rdrow_end          : in    std_logic := 'U';
          Sdram_ctl_v2_0_SD_rdEN_noact   : in    std_logic := 'U'
        );
  end component;

  component Main_ctl4SD
    port( intData2acc_RNIPB46                 : out   std_logic_vector(71 to 71);
          intData2acc_RNIFHV6                 : out   std_logic_vector(4 to 4);
          intData2acc_RNIEDV6                 : out   std_logic_vector(3 to 3);
          intData2acc_RNIITV6                 : out   std_logic_vector(7 to 7);
          intData2acc_RNIHPV6                 : out   std_logic_vector(6 to 6);
          intData2acc_RNIGLV6                 : out   std_logic_vector(5 to 5);
          intData2acc_RNI6J36                 : out   std_logic_vector(10 to 10);
          intData2acc_RNIK507                 : out   std_logic_vector(9 to 9);
          intData2acc_RNIJ107                 : out   std_logic_vector(8 to 8);
          intData2acc_RNI9J36                 : out   std_logic_vector(13 to 13);
          intData2acc_RNI8J36                 : out   std_logic_vector(12 to 12);
          intData2acc_RNI7J36                 : out   std_logic_vector(11 to 11);
          intData2acc_RNICJ36                 : out   std_logic_vector(16 to 16);
          intData2acc_RNIBJ36                 : out   std_logic_vector(15 to 15);
          intData2acc_RNIAJ36                 : out   std_logic_vector(14 to 14);
          intData2acc_RNIDJ36                 : out   std_logic_vector(17 to 17);
          intData2acc_RNIBN36                 : out   std_logic_vector(22 to 22);
          intData2acc_RNIAN36                 : out   std_logic_vector(21 to 21);
          intData2acc_RNIEN36                 : out   std_logic_vector(25 to 25);
          intData2acc_RNIDN36                 : out   std_logic_vector(24 to 24);
          intData2acc_RNITJS7                 : out   std_logic_vector(23 to 23);
          intData2acc_RNI2KS7                 : out   std_logic_vector(28 to 28);
          intData2acc_RNI1KS7                 : out   std_logic_vector(27 to 27);
          intData2acc_RNI0KS7                 : out   std_logic_vector(26 to 26);
          intData2acc_RNI4JV9                 : out   std_logic_vector(31 to 31);
          intData2acc_RNI3JV9                 : out   std_logic_vector(30 to 30);
          intData2acc_RNI9FV9                 : out   std_logic_vector(29 to 29);
          intData2acc_RNI5JV9                 : out   std_logic_vector(32 to 32);
          intData2acc_RNI8JV9                 : out   std_logic_vector(35 to 35);
          intData2acc_RNI6NV9                 : out   std_logic_vector(40 to 40);
          intData2acc_RNICJV9                 : out   std_logic_vector(39 to 39);
          intData2acc_RNIBJV9                 : out   std_logic_vector(38 to 38);
          intData2acc_RNI9NV9                 : out   std_logic_vector(43 to 43);
          intData2acc_RNI8NV9                 : out   std_logic_vector(42 to 42);
          intData2acc_RNI7NV9                 : out   std_logic_vector(41 to 41);
          intData2acc_RNICNV9                 : out   std_logic_vector(46 to 46);
          intData2acc_RNIBNV9                 : out   std_logic_vector(45 to 45);
          intData2acc_RNIANV9                 : out   std_logic_vector(44 to 44);
          intData2acc_RNIFNV9                 : out   std_logic_vector(49 to 49);
          intData2acc_RNIENV9                 : out   std_logic_vector(48 to 48);
          intData2acc_RNIDNV9                 : out   std_logic_vector(47 to 47);
          intData2acc_RNI9RV9                 : out   std_logic_vector(51 to 51);
          intData2acc_RNI8RV9                 : out   std_logic_vector(50 to 50);
          intData2acc_RNIERV9                 : out   std_logic_vector(57 to 57);
          intData2acc_RNIDRV9                 : out   std_logic_vector(56 to 56);
          intData2acc_RNIBVV9                 : out   std_logic_vector(61 to 61);
          intData2acc_RNIAVV9                 : out   std_logic_vector(60 to 60);
          intData2acc_RNIGRV9                 : out   std_logic_vector(59 downto 58);
          intData2acc_RNIEVV9                 : out   std_logic_vector(64 to 64);
          intData2acc_RNIDVV9                 : out   std_logic_vector(63 to 63);
          intData2acc_RNICVV9                 : out   std_logic_vector(62 to 62);
          intData2acc_RNIHVV9                 : out   std_logic_vector(67 to 67);
          intData2acc_RNIGVV9                 : out   std_logic_vector(66 to 66);
          intData2acc_RNIFVV9                 : out   std_logic_vector(65 to 65);
          intData2acc_RNID30A                 : out   std_logic_vector(70 to 70);
          intData2acc_RNIVOQA                 : out   std_logic_vector(0 to 0);
          intData2acc_RNI2BV9                 : out   std_logic_vector(18 to 18);
          intData2acc_RNI6JV9_0               : out   std_logic;
          intData2acc_RNI6JV9_3               : out   std_logic;
          intData2acc_RNI0TQA                 : out   std_logic_vector(1 to 1);
          intData2acc_RNI3BV9                 : out   std_logic_vector(19 to 19);
          intData2acc_RNI7JV9_0               : out   std_logic;
          intData2acc_RNI7JV9_3               : out   std_logic;
          intData2acc_RNI11RA                 : out   std_logic_vector(2 to 2);
          intData2acc_RNITEV9                 : out   std_logic_vector(20 to 20);
          pr_state_ns                         : in    std_logic_vector(8 to 8) := (others => 'U');
          intData2acc_RNIARV9                 : out   std_logic_vector(54 to 54);
          intData2acc_RNIBRV9_0               : out   std_logic;
          intData2acc_RNIBRV9_1               : out   std_logic;
          intData2acc_RNIBRV9_3               : out   std_logic;
          Main_ctl4SD_0_ByteRdEn              : out   std_logic;
          CMOS_DrvX_0_LVDSen_1                : in    std_logic := 'U';
          CMOS_DrvX_0_LVDSen_2                : in    std_logic := 'U';
          Main_ctl4SD_0_Fifo_wr               : out   std_logic;
          Main_ctl4SD_0_fifo_rd               : out   std_logic;
          \Z\\Fifo_rd_0_Q_[71]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[70]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[69]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[68]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[67]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[66]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[65]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[64]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[63]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[62]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[61]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[60]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[59]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[58]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[57]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[56]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[55]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[54]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[53]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[52]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[51]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[50]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[49]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[48]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[47]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[46]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[45]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[44]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[43]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[42]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[41]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[40]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[39]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[38]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[37]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[36]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[35]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[34]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[33]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[32]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[31]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[30]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[29]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[28]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[27]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[26]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[25]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[24]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[23]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[22]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[21]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[20]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[19]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[18]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[17]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[16]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[15]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[14]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[13]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[12]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[11]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[10]\\\             : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[9]\\\              : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[8]\\\              : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[7]\\\              : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[6]\\\              : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[5]\\\              : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[4]\\\              : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[3]\\\              : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[2]\\\              : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[1]\\\              : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[0]\\\              : in    std_logic := 'U';
          CMOS_DrvX_0_SDramEn_2               : in    std_logic := 'U';
          CMOS_DrvX_0_SDramEn_1               : in    std_logic := 'U';
          CMOS_DrvX_0_SDramEn                 : in    std_logic := 'U';
          CMOS_DrvX_0_SDramEn_5               : in    std_logic := 'U';
          CMOS_DrvX_0_SDramEn_4               : in    std_logic := 'U';
          CMOS_DrvX_0_SDramEn_3               : in    std_logic := 'U';
          \Z\\Main_ctl4SD_0_Data2Fifo_[71]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[70]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[69]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[68]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[67]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[66]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[65]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[64]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[63]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[62]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[61]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[60]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[59]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[58]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[57]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[56]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[55]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[54]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[53]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[52]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[51]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[50]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[49]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[48]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[47]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[46]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[45]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[44]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[43]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[42]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[41]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[40]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[39]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[38]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[37]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[36]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[35]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[34]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[33]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[32]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[31]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[30]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[29]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[28]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[27]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[26]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[25]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[24]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[23]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[22]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[21]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[20]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[19]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[18]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[17]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[16]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[15]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[14]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[13]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[12]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[11]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[10]\\\ : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[9]\\\  : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[8]\\\  : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[7]\\\  : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[6]\\\  : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[5]\\\  : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[4]\\\  : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[3]\\\  : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[2]\\\  : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[1]\\\  : out   std_logic;
          \Z\\Main_ctl4SD_0_Data2Fifo_[0]\\\  : out   std_logic;
          Main_ctl4SD_0_fifo_rst_n            : out   std_logic;
          FrameMk_0_LVDS_ok                   : in    std_logic := 'U';
          CMOS_DrvX_0_SDramEn_0               : in    std_logic := 'U';
          LVDS_enReg                          : in    std_logic := 'U';
          un6_sdramenreg                      : out   std_logic;
          CMOS_DrvX_0_AdcEn                   : in    std_logic := 'U';
          N_6                                 : out   std_logic;
          N_4                                 : out   std_logic;
          \Z\\My_adder0_0_Sum_[3]\\\          : in    std_logic := 'U';
          \Z\\My_adder0_0_Sum_[2]\\\          : in    std_logic := 'U';
          \Z\\My_adder0_0_Sum_[1]\\\          : in    std_logic := 'U';
          \Z\\My_adder0_0_Sum_[0]\\\          : in    std_logic := 'U';
          \Z\\My_adder0_0_Sum_[7]\\\          : in    std_logic := 'U';
          \Z\\My_adder0_0_Sum_[6]\\\          : in    std_logic := 'U';
          \Z\\My_adder0_0_Sum_[5]\\\          : in    std_logic := 'U';
          \Z\\My_adder0_0_Sum_[4]\\\          : in    std_logic := 'U';
          \Z\\My_adder0_0_Sum_[11]\\\         : in    std_logic := 'U';
          \Z\\My_adder0_0_Sum_[10]\\\         : in    std_logic := 'U';
          \Z\\My_adder0_0_Sum_[9]\\\          : in    std_logic := 'U';
          \Z\\My_adder0_0_Sum_[8]\\\          : in    std_logic := 'U';
          \Z\\My_adder0_0_Sum_[15]\\\         : in    std_logic := 'U';
          \Z\\My_adder0_0_Sum_[14]\\\         : in    std_logic := 'U';
          \Z\\My_adder0_0_Sum_[13]\\\         : in    std_logic := 'U';
          \Z\\My_adder0_0_Sum_[12]\\\         : in    std_logic := 'U';
          \Z\\My_adder0_2_Sum_[1]\\\          : in    std_logic := 'U';
          \Z\\My_adder0_2_Sum_[0]\\\          : in    std_logic := 'U';
          \Z\\My_adder0_1_Sum_[8]\\\          : in    std_logic := 'U';
          \Z\\My_adder0_0_Sum_[16]\\\         : in    std_logic := 'U';
          \Z\\My_adder0_2_Sum_[3]\\\          : in    std_logic := 'U';
          \Z\\My_adder0_2_Sum_[2]\\\          : in    std_logic := 'U';
          \Z\\My_adder0_1_Sum_[9]\\\          : in    std_logic := 'U';
          \Z\\My_adder0_0_Sum_[17]\\\         : in    std_logic := 'U';
          \Z\\My_adder0_2_Sum_[5]\\\          : in    std_logic := 'U';
          \Z\\My_adder0_2_Sum_[4]\\\          : in    std_logic := 'U';
          \Z\\My_adder0_1_Sum_[10]\\\         : in    std_logic := 'U';
          \Z\\My_adder0_1_Sum_[0]\\\          : in    std_logic := 'U';
          \Z\\My_adder0_2_Sum_[7]\\\          : in    std_logic := 'U';
          \Z\\My_adder0_2_Sum_[6]\\\          : in    std_logic := 'U';
          \Z\\My_adder0_1_Sum_[11]\\\         : in    std_logic := 'U';
          \Z\\My_adder0_1_Sum_[1]\\\          : in    std_logic := 'U';
          \Z\\My_adder0_2_Sum_[9]\\\          : in    std_logic := 'U';
          \Z\\My_adder0_2_Sum_[8]\\\          : in    std_logic := 'U';
          \Z\\My_adder0_1_Sum_[12]\\\         : in    std_logic := 'U';
          \Z\\My_adder0_1_Sum_[2]\\\          : in    std_logic := 'U';
          \Z\\My_adder0_2_Sum_[11]\\\         : in    std_logic := 'U';
          \Z\\My_adder0_2_Sum_[10]\\\         : in    std_logic := 'U';
          \Z\\My_adder0_1_Sum_[13]\\\         : in    std_logic := 'U';
          \Z\\My_adder0_1_Sum_[3]\\\          : in    std_logic := 'U';
          \Z\\My_adder0_2_Sum_[13]\\\         : in    std_logic := 'U';
          \Z\\My_adder0_2_Sum_[12]\\\         : in    std_logic := 'U';
          \Z\\My_adder0_1_Sum_[14]\\\         : in    std_logic := 'U';
          \Z\\My_adder0_1_Sum_[4]\\\          : in    std_logic := 'U';
          \Z\\My_adder0_2_Sum_[15]\\\         : in    std_logic := 'U';
          \Z\\My_adder0_2_Sum_[14]\\\         : in    std_logic := 'U';
          \Z\\My_adder0_1_Sum_[15]\\\         : in    std_logic := 'U';
          \Z\\My_adder0_1_Sum_[5]\\\          : in    std_logic := 'U';
          \Z\\My_adder0_2_Sum_[17]\\\         : in    std_logic := 'U';
          \Z\\My_adder0_2_Sum_[16]\\\         : in    std_logic := 'U';
          \Z\\My_adder0_1_Sum_[16]\\\         : in    std_logic := 'U';
          \Z\\My_adder0_1_Sum_[6]\\\          : in    std_logic := 'U';
          \Z\\My_adder0_3_Sum_[1]\\\          : in    std_logic := 'U';
          \Z\\My_adder0_3_Sum_[0]\\\          : in    std_logic := 'U';
          \Z\\My_adder0_1_Sum_[17]\\\         : in    std_logic := 'U';
          \Z\\My_adder0_1_Sum_[7]\\\          : in    std_logic := 'U';
          \Z\\My_adder0_3_Sum_[5]\\\          : in    std_logic := 'U';
          \Z\\My_adder0_3_Sum_[4]\\\          : in    std_logic := 'U';
          \Z\\My_adder0_3_Sum_[3]\\\          : in    std_logic := 'U';
          \Z\\My_adder0_3_Sum_[2]\\\          : in    std_logic := 'U';
          \Z\\My_adder0_3_Sum_[9]\\\          : in    std_logic := 'U';
          \Z\\My_adder0_3_Sum_[8]\\\          : in    std_logic := 'U';
          \Z\\My_adder0_3_Sum_[7]\\\          : in    std_logic := 'U';
          \Z\\My_adder0_3_Sum_[6]\\\          : in    std_logic := 'U';
          \Z\\My_adder0_3_Sum_[13]\\\         : in    std_logic := 'U';
          \Z\\My_adder0_3_Sum_[12]\\\         : in    std_logic := 'U';
          \Z\\My_adder0_3_Sum_[11]\\\         : in    std_logic := 'U';
          \Z\\My_adder0_3_Sum_[10]\\\         : in    std_logic := 'U';
          \Z\\My_adder0_3_Sum_[17]\\\         : in    std_logic := 'U';
          \Z\\My_adder0_3_Sum_[16]\\\         : in    std_logic := 'U';
          \Z\\My_adder0_3_Sum_[15]\\\         : in    std_logic := 'U';
          \Z\\My_adder0_3_Sum_[14]\\\         : in    std_logic := 'U';
          FrameMk_0_LVDS_ok_i                 : in    std_logic := 'U';
          Main_ctl4SD_0_fifo_rst_n_0          : out   std_logic;
          Main_ctl4SD_0_fifo_rst_n_1          : out   std_logic;
          Main_ctl4SD_0_fifo_rst_n_2          : out   std_logic;
          Main_ctl4SD_0_fifo_rst_n_3          : out   std_logic;
          Main_ctl4SD_0_fifo_rst_n_4          : out   std_logic;
          Main_ctl4SD_0_fifo_rst_n_5          : out   std_logic;
          PLL_Test1_0_SysRst_O                : in    std_logic := 'U';
          PLL_Test1_0_Sys_66M_Clk             : in    std_logic := 'U';
          Main_ctl4SD_0_fifo_rst_n_6          : out   std_logic
        );
  end component;

  component Fifo_rd_1
    port( \Z\\Fifo_rd_0_Q_[27]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[23]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[69]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[1]\\\               : out   std_logic;
          \Z\\Fifo_rd_0_Q_[67]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[4]\\\               : out   std_logic;
          \Z\\Fifo_rd_0_Q_[63]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[7]\\\               : out   std_logic;
          \Z\\Fifo_rd_0_Q_[56]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[25]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[24]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[48]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[65]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[64]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[51]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[38]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[71]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[50]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[70]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[18]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[6]\\\               : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[71]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[70]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[69]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[68]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[67]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[66]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[65]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[64]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[63]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[62]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[61]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[60]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[59]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[58]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[57]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[56]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[55]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[54]\\\ : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[46]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[52]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[36]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[59]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[0]\\\               : out   std_logic;
          \Z\\Fifo_rd_0_Q_[16]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[57]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[41]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[53]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[40]\\\              : out   std_logic;
          Main_ctl4SD_0_fifo_rd                : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[31]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[28]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[30]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[42]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[11]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[10]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[55]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[68]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[54]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[49]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[9]\\\               : out   std_logic;
          \Z\\Fifo_rd_0_Q_[5]\\\               : out   std_logic;
          Fifo_rd_0_AFULL                      : out   std_logic;
          \Z\\Fifo_rd_0_Q_[32]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[47]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[43]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[12]\\\              : out   std_logic;
          Sdram_cmd_0_RFifo_we                 : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[26]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[39]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[19]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[37]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[3]\\\               : out   std_logic;
          \Z\\Fifo_rd_0_Q_[33]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[66]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[17]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[13]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[45]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[44]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[21]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[2]\\\               : out   std_logic;
          \Z\\Fifo_rd_0_Q_[20]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[61]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[35]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[34]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[60]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[15]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[14]\\\              : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[35]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[34]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[33]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[32]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[31]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[30]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[29]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[28]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[27]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[26]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[25]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[24]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[23]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[22]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[21]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[20]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[19]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[18]\\\ : in    std_logic := 'U';
          Main_ctl4SD_0_fifo_rst_n_0           : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[22]\\\              : out   std_logic;
          \Z\\Fifo_rd_0_Q_[8]\\\               : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[53]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[52]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[51]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[50]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[49]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[48]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[47]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[46]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[45]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[44]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[43]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[42]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[41]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[40]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[39]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[38]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[37]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[36]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[17]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[16]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[15]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[14]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[13]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[12]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[11]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[10]\\\ : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[9]\\\  : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[8]\\\  : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[7]\\\  : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[6]\\\  : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[5]\\\  : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[4]\\\  : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[3]\\\  : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[2]\\\  : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[1]\\\  : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[0]\\\  : in    std_logic := 'U';
          Fifo_rd_1_VCC                        : in    std_logic := 'U';
          Main_ctl4SD_0_fifo_rst_n_3           : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[62]\\\              : out   std_logic;
          Main_ctl4SD_0_fifo_rst_n_1           : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[29]\\\              : out   std_logic;
          Main_ctl4SD_0_fifo_rst_n_2           : in    std_logic := 'U';
          PLL_Test1_0_Sys_66M_Clk              : in    std_logic := 'U';
          \Z\\Fifo_rd_0_Q_[58]\\\              : out   std_logic;
          Fifo_rd_1_GND                        : in    std_logic := 'U'
        );
  end component;

  component Sdram_data
    port( Sd_DQ_in                             : in    std_logic_vector(71 downto 0) := (others => 'U');
          \Z\\Sdram_data_0_Sys_dataOut_[71]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[70]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[69]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[68]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[67]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[66]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[65]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[64]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[63]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[62]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[61]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[60]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[59]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[58]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[57]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[56]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[55]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[54]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[53]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[52]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[51]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[50]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[49]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[48]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[47]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[46]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[45]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[44]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[43]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[42]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[41]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[40]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[39]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[38]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[37]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[36]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[35]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[34]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[33]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[32]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[31]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[30]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[29]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[28]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[27]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[26]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[25]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[24]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[23]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[22]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[21]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[20]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[19]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[18]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[17]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[16]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[15]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[14]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[13]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[12]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[11]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[10]\\\ : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[9]\\\  : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[8]\\\  : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[7]\\\  : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[6]\\\  : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[5]\\\  : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[4]\\\  : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[3]\\\  : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[2]\\\  : out   std_logic;
          \Z\\Sdram_data_0_Sys_dataOut_[1]\\\  : out   std_logic;
          PLL_Test1_0_SysRst_O                 : in    std_logic := 'U';
          PLL_Test1_0_Sys_66M_Clk              : in    std_logic := 'U';
          \Z\\Sdram_data_0_Sys_dataOut_[0]\\\  : out   std_logic;
          \Z\\SDram_rd_0_rd_state_[1]\\\       : in    std_logic := 'U';
          \Z\\SDram_rd_0_rd_state_[2]\\\       : in    std_logic := 'U';
          \Z\\SDram_rd_0_rd_state_[0]\\\       : in    std_logic := 'U'
        );
  end component;

  component adc_muxtmp_test
    port( PLL_Test1_0_SysRst_O                        : in    std_logic := 'U';
          PLL_Test1_0_Sys_66M_Clk                     : in    std_logic := 'U';
          CMOS_DrvX_0_AdcEn                           : in    std_logic := 'U';
          \Z\\adc_muxtmp_test_0_DataOut41to28_[29]\\\ : out   std_logic;
          \Z\\adc_muxtmp_test_0_DataOut27to14_[14]\\\ : out   std_logic;
          \Z\\adc_muxtmp_test_0_DataOut55to42_[43]\\\ : out   std_logic
        );
  end component;

  component PLL_Test1
    port( PLL_Test1_0_ADC_66M_Clk : out   std_logic;
          PLL_Test1_0_Sdram_clk   : out   std_logic;
          ExterCLk_c              : in    std_logic := 'U';
          PLL_Test1_GND           : in    std_logic := 'U';
          PLL_Test1_0_SysRst_O    : out   std_logic;
          PLL_Test1_VCC           : in    std_logic := 'U';
          PLL_Test1_0_Sys_66M_Clk : out   std_logic
        );
  end component;

  component Sdram_ctl_v2
    port( SD_cke_c_c                   : out   std_logic_vector(0 to 0);
          pr_state_ns_3                : out   std_logic;
          Sdram_ini_0_Sd_iniOK_i       : in    std_logic := 'U';
          Sdram_ctl_v2_0_SD_iniEn      : out   std_logic;
          Sdram_ctl_v2_0_SD_RefEn      : out   std_logic;
          Sdram_ctl_v2_0_SD_rdEN_noact : out   std_logic;
          PLL_Test1_0_SysRst_O         : in    std_logic := 'U';
          PLL_Test1_0_Sys_66M_Clk      : in    std_logic := 'U';
          Sdram_ctl_v2_0_SD_pdEN       : out   std_logic;
          Fifo_wr_0_AFULL              : in    std_logic := 'U';
          SDRAM_wr_0_SD_WrOK           : in    std_logic := 'U';
          ref_ok_2                     : in    std_logic := 'U';
          ref_ok_1                     : in    std_logic := 'U';
          CMOS_DrvX_0_LVDSen_2         : in    std_logic := 'U';
          CMOS_DrvX_0_SDramEn_0        : in    std_logic := 'U';
          Sdram_ini_0_Sd_iniOK         : in    std_logic := 'U';
          Fifo_rd_0_AFULL              : in    std_logic := 'U';
          CMOS_DrvX_0_LVDSen_1         : in    std_logic := 'U';
          SDram_rd_0_SD_RdOK           : in    std_logic := 'U';
          Sdram_ctl_v2_0_SD_rdEn       : out   std_logic;
          Sdram_ctl_v2_0_SD_rdEn_i     : out   std_logic;
          Sdram_ctl_v2_0_SD_wrEn       : out   std_logic;
          Sdram_ctl_v2_0_SD_wrEn_i     : out   std_logic
        );
  end component;

  component My_adder0_2
    port( intData2acc_RNI2KS7                         : in    std_logic_vector(28 to 28) := (others => 'U');
          intData2acc_RNI1KS7                         : in    std_logic_vector(27 to 27) := (others => 'U');
          intData2acc_RNI6JV9                         : in    std_logic_vector(33 to 33) := (others => 'U');
          intData2acc_RNI2BV9                         : in    std_logic_vector(18 to 18) := (others => 'U');
          intData2acc_RNI3BV9                         : in    std_logic_vector(19 to 19) := (others => 'U');
          intData2acc_RNIBN36                         : in    std_logic_vector(22 to 22) := (others => 'U');
          intData2acc_RNI3JV9                         : in    std_logic_vector(30 to 30) := (others => 'U');
          intData2acc_RNI5JV9                         : in    std_logic_vector(32 to 32) := (others => 'U');
          intData2acc_RNITEV9                         : in    std_logic_vector(20 to 20) := (others => 'U');
          intData2acc_RNIAN36                         : in    std_logic_vector(21 to 21) := (others => 'U');
          intData2acc_RNI4JV9                         : in    std_logic_vector(31 to 31) := (others => 'U');
          intData2acc_RNIDN36                         : in    std_logic_vector(24 to 24) := (others => 'U');
          intData2acc_RNIEN36                         : in    std_logic_vector(25 to 25) := (others => 'U');
          intData2acc_RNI9FV9                         : in    std_logic_vector(29 to 29) := (others => 'U');
          intData2acc_RNI8JV9                         : in    std_logic_vector(35 to 35) := (others => 'U');
          intData2acc_RNITJS7                         : in    std_logic_vector(23 to 23) := (others => 'U');
          intData2acc_RNI0KS7                         : in    std_logic_vector(26 to 26) := (others => 'U');
          intData2acc_RNI7JV9                         : in    std_logic_vector(34 to 34) := (others => 'U');
          \Z\\My_adder0_1_Sum_[15]\\\                 : out   std_logic;
          \Z\\My_adder0_1_Sum_[12]\\\                 : out   std_logic;
          \Z\\My_adder0_1_Sum_[6]\\\                  : out   std_logic;
          \Z\\My_adder0_1_Sum_[10]\\\                 : out   std_logic;
          \Z\\My_adder0_1_Sum_[9]\\\                  : out   std_logic;
          \Z\\My_adder0_1_Sum_[7]\\\                  : out   std_logic;
          \Z\\My_adder0_1_Sum_[11]\\\                 : out   std_logic;
          \Z\\My_adder0_1_Sum_[1]\\\                  : out   std_logic;
          \Z\\My_adder0_1_Sum_[3]\\\                  : out   std_logic;
          \Z\\My_adder0_1_Sum_[13]\\\                 : out   std_logic;
          \Z\\adc_muxtmp_test_0_DataOut27to14_[14]\\\ : in    std_logic := 'U';
          \Z\\My_adder0_1_Sum_[0]\\\                  : out   std_logic;
          \Z\\My_adder0_1_Sum_[8]\\\                  : out   std_logic;
          \Z\\My_adder0_1_Sum_[14]\\\                 : out   std_logic;
          \Z\\My_adder0_1_Sum_[2]\\\                  : out   std_logic;
          \Z\\My_adder0_1_Sum_[4]\\\                  : out   std_logic;
          \Z\\My_adder0_1_Sum_[5]\\\                  : out   std_logic;
          \Z\\My_adder0_1_Sum_[17]\\\                 : out   std_logic;
          My_adder0_2_GND                             : in    std_logic := 'U';
          \Z\\My_adder0_1_Sum_[16]\\\                 : out   std_logic
        );
  end component;

    signal \My_adder0_2_Sum_[0]\, \My_adder0_2_Sum_[1]\, 
        \My_adder0_2_Sum_[2]\, \My_adder0_2_Sum_[3]\, 
        \My_adder0_2_Sum_[4]\, \My_adder0_2_Sum_[5]\, 
        \My_adder0_2_Sum_[6]\, \My_adder0_2_Sum_[7]\, 
        \My_adder0_2_Sum_[8]\, \My_adder0_2_Sum_[9]\, 
        \My_adder0_2_Sum_[10]\, \My_adder0_2_Sum_[11]\, 
        \My_adder0_2_Sum_[12]\, \My_adder0_2_Sum_[13]\, 
        \My_adder0_2_Sum_[14]\, \My_adder0_2_Sum_[15]\, 
        \My_adder0_2_Sum_[16]\, \My_adder0_2_Sum_[17]\, 
        \Fifo_wr_0_Q_[0]\, \Fifo_wr_0_Q_[1]\, \Fifo_wr_0_Q_[2]\, 
        \Fifo_wr_0_Q_[3]\, \Fifo_wr_0_Q_[4]\, \Fifo_wr_0_Q_[5]\, 
        \Fifo_wr_0_Q_[6]\, \Fifo_wr_0_Q_[7]\, \Fifo_wr_0_Q_[8]\, 
        \Fifo_wr_0_Q_[9]\, \Fifo_wr_0_Q_[10]\, \Fifo_wr_0_Q_[11]\, 
        \Fifo_wr_0_Q_[12]\, \Fifo_wr_0_Q_[13]\, 
        \Fifo_wr_0_Q_[14]\, \Fifo_wr_0_Q_[15]\, 
        \Fifo_wr_0_Q_[16]\, \Fifo_wr_0_Q_[17]\, 
        \Fifo_wr_0_Q_[18]\, \Fifo_wr_0_Q_[19]\, 
        \Fifo_wr_0_Q_[20]\, \Fifo_wr_0_Q_[21]\, 
        \Fifo_wr_0_Q_[22]\, \Fifo_wr_0_Q_[23]\, 
        \Fifo_wr_0_Q_[24]\, \Fifo_wr_0_Q_[25]\, 
        \Fifo_wr_0_Q_[26]\, \Fifo_wr_0_Q_[27]\, 
        \Fifo_wr_0_Q_[28]\, \Fifo_wr_0_Q_[29]\, 
        \Fifo_wr_0_Q_[30]\, \Fifo_wr_0_Q_[31]\, 
        \Fifo_wr_0_Q_[32]\, \Fifo_wr_0_Q_[33]\, 
        \Fifo_wr_0_Q_[34]\, \Fifo_wr_0_Q_[35]\, 
        \Fifo_wr_0_Q_[36]\, \Fifo_wr_0_Q_[37]\, 
        \Fifo_wr_0_Q_[38]\, \Fifo_wr_0_Q_[39]\, 
        \Fifo_wr_0_Q_[40]\, \Fifo_wr_0_Q_[41]\, 
        \Fifo_wr_0_Q_[42]\, \Fifo_wr_0_Q_[43]\, 
        \Fifo_wr_0_Q_[44]\, \Fifo_wr_0_Q_[45]\, 
        \Fifo_wr_0_Q_[46]\, \Fifo_wr_0_Q_[47]\, 
        \Fifo_wr_0_Q_[48]\, \Fifo_wr_0_Q_[49]\, 
        \Fifo_wr_0_Q_[50]\, \Fifo_wr_0_Q_[51]\, 
        \Fifo_wr_0_Q_[52]\, \Fifo_wr_0_Q_[53]\, 
        \Fifo_wr_0_Q_[54]\, \Fifo_wr_0_Q_[55]\, 
        \Fifo_wr_0_Q_[56]\, \Fifo_wr_0_Q_[57]\, 
        \Fifo_wr_0_Q_[58]\, \Fifo_wr_0_Q_[59]\, 
        \Fifo_wr_0_Q_[60]\, \Fifo_wr_0_Q_[61]\, 
        \Fifo_wr_0_Q_[62]\, \Fifo_wr_0_Q_[63]\, 
        \Fifo_wr_0_Q_[64]\, \Fifo_wr_0_Q_[65]\, 
        \Fifo_wr_0_Q_[66]\, \Fifo_wr_0_Q_[67]\, 
        \Fifo_wr_0_Q_[68]\, \Fifo_wr_0_Q_[69]\, 
        \Fifo_wr_0_Q_[70]\, \Fifo_wr_0_Q_[71]\, 
        Main_ctl4SD_0_Fifo_wr, Sdram_cmd_0_WFifo_re, 
        PLL_Test1_0_Sys_66M_Clk, Main_ctl4SD_0_fifo_rst_n, 
        Fifo_wr_0_AFULL, PLL_Test1_0_SysRst_O, 
        \adc_muxtmp_test_0_DataOut27to14_[14]\, 
        \adc_muxtmp_test_0_DataOut41to28_[29]\, 
        \adc_muxtmp_test_0_DataOut55to42_[43]\, 
        Sdram_ctl_v2_0_SD_iniEn, Sdram_ini_0_Sd_iniOK, 
        \Sdram_ini_0_ini_state_[0]\, \Sdram_ini_0_ini_state_[1]\, 
        \Sdram_ini_0_ini_state_[2]\, \My_adder0_3_Sum_[0]\, 
        \My_adder0_3_Sum_[1]\, \My_adder0_3_Sum_[2]\, 
        \My_adder0_3_Sum_[3]\, \My_adder0_3_Sum_[4]\, 
        \My_adder0_3_Sum_[5]\, \My_adder0_3_Sum_[6]\, 
        \My_adder0_3_Sum_[7]\, \My_adder0_3_Sum_[8]\, 
        \My_adder0_3_Sum_[9]\, \My_adder0_3_Sum_[10]\, 
        \My_adder0_3_Sum_[11]\, \My_adder0_3_Sum_[12]\, 
        \My_adder0_3_Sum_[13]\, \My_adder0_3_Sum_[14]\, 
        \My_adder0_3_Sum_[15]\, \My_adder0_3_Sum_[16]\, 
        \My_adder0_3_Sum_[17]\, PLL_Test1_0_ADC_66M_Clk, 
        PLL_Test1_0_Sdram_clk, \My_adder0_1_Sum_[0]\, 
        \My_adder0_1_Sum_[1]\, \My_adder0_1_Sum_[2]\, 
        \My_adder0_1_Sum_[3]\, \My_adder0_1_Sum_[4]\, 
        \My_adder0_1_Sum_[5]\, \My_adder0_1_Sum_[6]\, 
        \My_adder0_1_Sum_[7]\, \My_adder0_1_Sum_[8]\, 
        \My_adder0_1_Sum_[9]\, \My_adder0_1_Sum_[10]\, 
        \My_adder0_1_Sum_[11]\, \My_adder0_1_Sum_[12]\, 
        \My_adder0_1_Sum_[13]\, \My_adder0_1_Sum_[14]\, 
        \My_adder0_1_Sum_[15]\, \My_adder0_1_Sum_[16]\, 
        \My_adder0_1_Sum_[17]\, Sdram_ctl_v2_0_SD_RefEn, 
        CMOS_DrvX_0_LVDSen, Main_ctl4SD_0_ByteRdEn, 
        Sdram_cmd_0_SDoneFrameOk, FrameMk_0_LVDS_ok, 
        CMOS_DrvX_0_SDramEn, \Main_ctl4SD_0_Data2Fifo_[0]\, 
        \Main_ctl4SD_0_Data2Fifo_[1]\, 
        \Main_ctl4SD_0_Data2Fifo_[2]\, 
        \Main_ctl4SD_0_Data2Fifo_[3]\, 
        \Main_ctl4SD_0_Data2Fifo_[4]\, 
        \Main_ctl4SD_0_Data2Fifo_[5]\, 
        \Main_ctl4SD_0_Data2Fifo_[6]\, 
        \Main_ctl4SD_0_Data2Fifo_[7]\, 
        \Main_ctl4SD_0_Data2Fifo_[8]\, 
        \Main_ctl4SD_0_Data2Fifo_[9]\, 
        \Main_ctl4SD_0_Data2Fifo_[10]\, 
        \Main_ctl4SD_0_Data2Fifo_[11]\, 
        \Main_ctl4SD_0_Data2Fifo_[12]\, 
        \Main_ctl4SD_0_Data2Fifo_[13]\, 
        \Main_ctl4SD_0_Data2Fifo_[14]\, 
        \Main_ctl4SD_0_Data2Fifo_[15]\, 
        \Main_ctl4SD_0_Data2Fifo_[16]\, 
        \Main_ctl4SD_0_Data2Fifo_[17]\, 
        \Main_ctl4SD_0_Data2Fifo_[18]\, 
        \Main_ctl4SD_0_Data2Fifo_[19]\, 
        \Main_ctl4SD_0_Data2Fifo_[20]\, 
        \Main_ctl4SD_0_Data2Fifo_[21]\, 
        \Main_ctl4SD_0_Data2Fifo_[22]\, 
        \Main_ctl4SD_0_Data2Fifo_[23]\, 
        \Main_ctl4SD_0_Data2Fifo_[24]\, 
        \Main_ctl4SD_0_Data2Fifo_[25]\, 
        \Main_ctl4SD_0_Data2Fifo_[26]\, 
        \Main_ctl4SD_0_Data2Fifo_[27]\, 
        \Main_ctl4SD_0_Data2Fifo_[28]\, 
        \Main_ctl4SD_0_Data2Fifo_[29]\, 
        \Main_ctl4SD_0_Data2Fifo_[30]\, 
        \Main_ctl4SD_0_Data2Fifo_[31]\, 
        \Main_ctl4SD_0_Data2Fifo_[32]\, 
        \Main_ctl4SD_0_Data2Fifo_[33]\, 
        \Main_ctl4SD_0_Data2Fifo_[34]\, 
        \Main_ctl4SD_0_Data2Fifo_[35]\, 
        \Main_ctl4SD_0_Data2Fifo_[36]\, 
        \Main_ctl4SD_0_Data2Fifo_[37]\, 
        \Main_ctl4SD_0_Data2Fifo_[38]\, 
        \Main_ctl4SD_0_Data2Fifo_[39]\, 
        \Main_ctl4SD_0_Data2Fifo_[40]\, 
        \Main_ctl4SD_0_Data2Fifo_[41]\, 
        \Main_ctl4SD_0_Data2Fifo_[42]\, 
        \Main_ctl4SD_0_Data2Fifo_[43]\, 
        \Main_ctl4SD_0_Data2Fifo_[44]\, 
        \Main_ctl4SD_0_Data2Fifo_[45]\, 
        \Main_ctl4SD_0_Data2Fifo_[46]\, 
        \Main_ctl4SD_0_Data2Fifo_[47]\, 
        \Main_ctl4SD_0_Data2Fifo_[48]\, 
        \Main_ctl4SD_0_Data2Fifo_[49]\, 
        \Main_ctl4SD_0_Data2Fifo_[50]\, 
        \Main_ctl4SD_0_Data2Fifo_[51]\, 
        \Main_ctl4SD_0_Data2Fifo_[52]\, 
        \Main_ctl4SD_0_Data2Fifo_[53]\, 
        \Main_ctl4SD_0_Data2Fifo_[54]\, 
        \Main_ctl4SD_0_Data2Fifo_[55]\, 
        \Main_ctl4SD_0_Data2Fifo_[56]\, 
        \Main_ctl4SD_0_Data2Fifo_[57]\, 
        \Main_ctl4SD_0_Data2Fifo_[58]\, 
        \Main_ctl4SD_0_Data2Fifo_[59]\, 
        \Main_ctl4SD_0_Data2Fifo_[60]\, 
        \Main_ctl4SD_0_Data2Fifo_[61]\, 
        \Main_ctl4SD_0_Data2Fifo_[62]\, 
        \Main_ctl4SD_0_Data2Fifo_[63]\, 
        \Main_ctl4SD_0_Data2Fifo_[64]\, 
        \Main_ctl4SD_0_Data2Fifo_[65]\, 
        \Main_ctl4SD_0_Data2Fifo_[66]\, 
        \Main_ctl4SD_0_Data2Fifo_[67]\, 
        \Main_ctl4SD_0_Data2Fifo_[68]\, 
        \Main_ctl4SD_0_Data2Fifo_[69]\, 
        \Main_ctl4SD_0_Data2Fifo_[70]\, 
        \Main_ctl4SD_0_Data2Fifo_[71]\, Main_ctl4SD_0_fifo_rd, 
        \Fifo_rd_0_Q_[0]\, \Fifo_rd_0_Q_[1]\, \Fifo_rd_0_Q_[2]\, 
        \Fifo_rd_0_Q_[3]\, \Fifo_rd_0_Q_[4]\, \Fifo_rd_0_Q_[5]\, 
        \Fifo_rd_0_Q_[6]\, \Fifo_rd_0_Q_[7]\, \Fifo_rd_0_Q_[8]\, 
        \Fifo_rd_0_Q_[9]\, \Fifo_rd_0_Q_[10]\, \Fifo_rd_0_Q_[11]\, 
        \Fifo_rd_0_Q_[12]\, \Fifo_rd_0_Q_[13]\, 
        \Fifo_rd_0_Q_[14]\, \Fifo_rd_0_Q_[15]\, 
        \Fifo_rd_0_Q_[16]\, \Fifo_rd_0_Q_[17]\, 
        \Fifo_rd_0_Q_[18]\, \Fifo_rd_0_Q_[19]\, 
        \Fifo_rd_0_Q_[20]\, \Fifo_rd_0_Q_[21]\, 
        \Fifo_rd_0_Q_[22]\, \Fifo_rd_0_Q_[23]\, 
        \Fifo_rd_0_Q_[24]\, \Fifo_rd_0_Q_[25]\, 
        \Fifo_rd_0_Q_[26]\, \Fifo_rd_0_Q_[27]\, 
        \Fifo_rd_0_Q_[28]\, \Fifo_rd_0_Q_[29]\, 
        \Fifo_rd_0_Q_[30]\, \Fifo_rd_0_Q_[31]\, 
        \Fifo_rd_0_Q_[32]\, \Fifo_rd_0_Q_[33]\, 
        \Fifo_rd_0_Q_[34]\, \Fifo_rd_0_Q_[35]\, 
        \Fifo_rd_0_Q_[36]\, \Fifo_rd_0_Q_[37]\, 
        \Fifo_rd_0_Q_[38]\, \Fifo_rd_0_Q_[39]\, 
        \Fifo_rd_0_Q_[40]\, \Fifo_rd_0_Q_[41]\, 
        \Fifo_rd_0_Q_[42]\, \Fifo_rd_0_Q_[43]\, 
        \Fifo_rd_0_Q_[44]\, \Fifo_rd_0_Q_[45]\, 
        \Fifo_rd_0_Q_[46]\, \Fifo_rd_0_Q_[47]\, 
        \Fifo_rd_0_Q_[48]\, \Fifo_rd_0_Q_[49]\, 
        \Fifo_rd_0_Q_[50]\, \Fifo_rd_0_Q_[51]\, 
        \Fifo_rd_0_Q_[52]\, \Fifo_rd_0_Q_[53]\, 
        \Fifo_rd_0_Q_[54]\, \Fifo_rd_0_Q_[55]\, 
        \Fifo_rd_0_Q_[56]\, \Fifo_rd_0_Q_[57]\, 
        \Fifo_rd_0_Q_[58]\, \Fifo_rd_0_Q_[59]\, 
        \Fifo_rd_0_Q_[60]\, \Fifo_rd_0_Q_[61]\, 
        \Fifo_rd_0_Q_[62]\, \Fifo_rd_0_Q_[63]\, 
        \Fifo_rd_0_Q_[64]\, \Fifo_rd_0_Q_[65]\, 
        \Fifo_rd_0_Q_[66]\, \Fifo_rd_0_Q_[67]\, 
        \Fifo_rd_0_Q_[68]\, \Fifo_rd_0_Q_[69]\, 
        \Fifo_rd_0_Q_[70]\, \Fifo_rd_0_Q_[71]\, 
        Sdram_cmd_0_RFifo_we, Fifo_rd_0_AFULL, SDRAM_wr_0_SD_WrOK, 
        SDram_rd_0_SD_RdOK, Sdram_ctl_v2_0_SD_pdEN, 
        Sdram_ctl_v2_0_SD_wrEn, Sdram_ctl_v2_0_SD_rdEn, 
        Sdram_ctl_v2_0_SD_rdEN_noact, \SDRAM_Ref_0_Ref_state_[0]\, 
        \SDRAM_Ref_0_Ref_state_[1]\, \SDRAM_Ref_0_Ref_state_[2]\, 
        \Sdram_data_0_Sys_dataOut_[0]\, 
        \Sdram_data_0_Sys_dataOut_[1]\, 
        \Sdram_data_0_Sys_dataOut_[2]\, 
        \Sdram_data_0_Sys_dataOut_[3]\, 
        \Sdram_data_0_Sys_dataOut_[4]\, 
        \Sdram_data_0_Sys_dataOut_[5]\, 
        \Sdram_data_0_Sys_dataOut_[6]\, 
        \Sdram_data_0_Sys_dataOut_[7]\, 
        \Sdram_data_0_Sys_dataOut_[8]\, 
        \Sdram_data_0_Sys_dataOut_[9]\, 
        \Sdram_data_0_Sys_dataOut_[10]\, 
        \Sdram_data_0_Sys_dataOut_[11]\, 
        \Sdram_data_0_Sys_dataOut_[12]\, 
        \Sdram_data_0_Sys_dataOut_[13]\, 
        \Sdram_data_0_Sys_dataOut_[14]\, 
        \Sdram_data_0_Sys_dataOut_[15]\, 
        \Sdram_data_0_Sys_dataOut_[16]\, 
        \Sdram_data_0_Sys_dataOut_[17]\, 
        \Sdram_data_0_Sys_dataOut_[18]\, 
        \Sdram_data_0_Sys_dataOut_[19]\, 
        \Sdram_data_0_Sys_dataOut_[20]\, 
        \Sdram_data_0_Sys_dataOut_[21]\, 
        \Sdram_data_0_Sys_dataOut_[22]\, 
        \Sdram_data_0_Sys_dataOut_[23]\, 
        \Sdram_data_0_Sys_dataOut_[24]\, 
        \Sdram_data_0_Sys_dataOut_[25]\, 
        \Sdram_data_0_Sys_dataOut_[26]\, 
        \Sdram_data_0_Sys_dataOut_[27]\, 
        \Sdram_data_0_Sys_dataOut_[28]\, 
        \Sdram_data_0_Sys_dataOut_[29]\, 
        \Sdram_data_0_Sys_dataOut_[30]\, 
        \Sdram_data_0_Sys_dataOut_[31]\, 
        \Sdram_data_0_Sys_dataOut_[32]\, 
        \Sdram_data_0_Sys_dataOut_[33]\, 
        \Sdram_data_0_Sys_dataOut_[34]\, 
        \Sdram_data_0_Sys_dataOut_[35]\, 
        \Sdram_data_0_Sys_dataOut_[36]\, 
        \Sdram_data_0_Sys_dataOut_[37]\, 
        \Sdram_data_0_Sys_dataOut_[38]\, 
        \Sdram_data_0_Sys_dataOut_[39]\, 
        \Sdram_data_0_Sys_dataOut_[40]\, 
        \Sdram_data_0_Sys_dataOut_[41]\, 
        \Sdram_data_0_Sys_dataOut_[42]\, 
        \Sdram_data_0_Sys_dataOut_[43]\, 
        \Sdram_data_0_Sys_dataOut_[44]\, 
        \Sdram_data_0_Sys_dataOut_[45]\, 
        \Sdram_data_0_Sys_dataOut_[46]\, 
        \Sdram_data_0_Sys_dataOut_[47]\, 
        \Sdram_data_0_Sys_dataOut_[48]\, 
        \Sdram_data_0_Sys_dataOut_[49]\, 
        \Sdram_data_0_Sys_dataOut_[50]\, 
        \Sdram_data_0_Sys_dataOut_[51]\, 
        \Sdram_data_0_Sys_dataOut_[52]\, 
        \Sdram_data_0_Sys_dataOut_[53]\, 
        \Sdram_data_0_Sys_dataOut_[54]\, 
        \Sdram_data_0_Sys_dataOut_[55]\, 
        \Sdram_data_0_Sys_dataOut_[56]\, 
        \Sdram_data_0_Sys_dataOut_[57]\, 
        \Sdram_data_0_Sys_dataOut_[58]\, 
        \Sdram_data_0_Sys_dataOut_[59]\, 
        \Sdram_data_0_Sys_dataOut_[60]\, 
        \Sdram_data_0_Sys_dataOut_[61]\, 
        \Sdram_data_0_Sys_dataOut_[62]\, 
        \Sdram_data_0_Sys_dataOut_[63]\, 
        \Sdram_data_0_Sys_dataOut_[64]\, 
        \Sdram_data_0_Sys_dataOut_[65]\, 
        \Sdram_data_0_Sys_dataOut_[66]\, 
        \Sdram_data_0_Sys_dataOut_[67]\, 
        \Sdram_data_0_Sys_dataOut_[68]\, 
        \Sdram_data_0_Sys_dataOut_[69]\, 
        \Sdram_data_0_Sys_dataOut_[70]\, 
        \Sdram_data_0_Sys_dataOut_[71]\, Sdram_cmd_0_rdrow_end, 
        Sdram_cmd_0_wrrow_end, \SDram_rd_0_rd_state_[0]\, 
        \SDram_rd_0_rd_state_[1]\, \SDram_rd_0_rd_state_[2]\, 
        \SDRAM_wr_0_wr_state_[0]\, \SDRAM_wr_0_wr_state_[1]\, 
        \SDRAM_wr_0_wr_state_[2]\, \My_adder0_0_Sum_[0]\, 
        \My_adder0_0_Sum_[1]\, \My_adder0_0_Sum_[2]\, 
        \My_adder0_0_Sum_[3]\, \My_adder0_0_Sum_[4]\, 
        \My_adder0_0_Sum_[5]\, \My_adder0_0_Sum_[6]\, 
        \My_adder0_0_Sum_[7]\, \My_adder0_0_Sum_[8]\, 
        \My_adder0_0_Sum_[9]\, \My_adder0_0_Sum_[10]\, 
        \My_adder0_0_Sum_[11]\, \My_adder0_0_Sum_[12]\, 
        \My_adder0_0_Sum_[13]\, \My_adder0_0_Sum_[14]\, 
        \My_adder0_0_Sum_[15]\, \My_adder0_0_Sum_[16]\, 
        \My_adder0_0_Sum_[17]\, \VCC\, \Sdram_cmd_0.LVDS_enReg\, 
        \Sdram_cmd_0.N_264\, \SDRAM_Ref_0.ref_ok_1\, 
        \SDRAM_Ref_0.ref_ok_2\, \Sdram_ctl_v2_0.pr_state_ns[8]\, 
        \Main_ctl4SD_0.N_4\, \Main_ctl4SD_0.N_6\, 
        \intData2acc_RNID30A[70]\, \intData2acc_RNIFVV9[65]\, 
        \intData2acc_RNIGVV9[66]\, \intData2acc_RNIHVV9[67]\, 
        \intData2acc_RNICVV9[62]\, \intData2acc_RNIDVV9[63]\, 
        \intData2acc_RNIEVV9[64]\, \intData2acc_RNIGRV9[59]\, 
        \intData2acc_RNIAVV9[60]\, \intData2acc_RNIBVV9[61]\, 
        \intData2acc_RNIDRV9[56]\, \intData2acc_RNIERV9[57]\, 
        \intData2acc_RNIGRV9[58]\, \intData2acc_RNIBRV9[53]\, 
        \intData2acc_RNI8RV9[50]\, \intData2acc_RNI9RV9[51]\, 
        \intData2acc_RNIBRV9[52]\, \intData2acc_RNIDNV9[47]\, 
        \intData2acc_RNIENV9[48]\, \intData2acc_RNIFNV9[49]\, 
        \intData2acc_RNIANV9[44]\, \intData2acc_RNIBNV9[45]\, 
        \intData2acc_RNICNV9[46]\, \intData2acc_RNI7NV9[41]\, 
        \intData2acc_RNI8NV9[42]\, \intData2acc_RNI9NV9[43]\, 
        \intData2acc_RNIBJV9[38]\, \intData2acc_RNICJV9[39]\, 
        \intData2acc_RNI6NV9[40]\, \intData2acc_RNI8JV9[35]\, 
        \intData2acc_RNI5JV9[32]\, \intData2acc_RNI6JV9[33]\, 
        \intData2acc_RNI7JV9[34]\, \intData2acc_RNI9FV9[29]\, 
        \intData2acc_RNI3JV9[30]\, \intData2acc_RNI4JV9[31]\, 
        \intData2acc_RNI0KS7[26]\, \intData2acc_RNI1KS7[27]\, 
        \intData2acc_RNI2KS7[28]\, \intData2acc_RNITJS7[23]\, 
        \intData2acc_RNIDN36[24]\, \intData2acc_RNIEN36[25]\, 
        \intData2acc_RNIAN36[21]\, \intData2acc_RNIBN36[22]\, 
        \intData2acc_RNIDJ36[17]\, \intData2acc_RNIAJ36[14]\, 
        \intData2acc_RNIBJ36[15]\, \intData2acc_RNICJ36[16]\, 
        \intData2acc_RNI7J36[11]\, \intData2acc_RNI8J36[12]\, 
        \intData2acc_RNI9J36[13]\, \intData2acc_RNIJ107[8]\, 
        \intData2acc_RNIK507[9]\, \intData2acc_RNI6J36[10]\, 
        \intData2acc_RNIGLV6[5]\, \intData2acc_RNIHPV6[6]\, 
        \intData2acc_RNIITV6[7]\, \intData2acc_RNIEDV6[3]\, 
        \intData2acc_RNIFHV6[4]\, \intData2acc_RNIPB46[71]\, 
        \Sd_DQ_in[0]\, \Sd_DQ_in[1]\, \Sd_DQ_in[2]\, 
        \Sd_DQ_in[3]\, \Sd_DQ_in[4]\, \Sd_DQ_in[5]\, 
        \Sd_DQ_in[6]\, \Sd_DQ_in[7]\, \Sd_DQ_in[8]\, 
        \Sd_DQ_in[9]\, \Sd_DQ_in[10]\, \Sd_DQ_in[11]\, 
        \Sd_DQ_in[12]\, \Sd_DQ_in[13]\, \Sd_DQ_in[14]\, 
        \Sd_DQ_in[15]\, \Sd_DQ_in[16]\, \Sd_DQ_in[17]\, 
        \Sd_DQ_in[18]\, \Sd_DQ_in[19]\, \Sd_DQ_in[20]\, 
        \Sd_DQ_in[21]\, \Sd_DQ_in[22]\, \Sd_DQ_in[23]\, 
        \Sd_DQ_in[24]\, \Sd_DQ_in[25]\, \Sd_DQ_in[26]\, 
        \Sd_DQ_in[27]\, \Sd_DQ_in[28]\, \Sd_DQ_in[29]\, 
        \Sd_DQ_in[30]\, \Sd_DQ_in[31]\, \Sd_DQ_in[32]\, 
        \Sd_DQ_in[33]\, \Sd_DQ_in[34]\, \Sd_DQ_in[35]\, 
        \Sd_DQ_in[36]\, \Sd_DQ_in[37]\, \Sd_DQ_in[38]\, 
        \Sd_DQ_in[39]\, \Sd_DQ_in[40]\, \Sd_DQ_in[41]\, 
        \Sd_DQ_in[42]\, \Sd_DQ_in[43]\, \Sd_DQ_in[44]\, 
        \Sd_DQ_in[45]\, \Sd_DQ_in[46]\, \Sd_DQ_in[47]\, 
        \Sd_DQ_in[48]\, \Sd_DQ_in[49]\, \Sd_DQ_in[50]\, 
        \Sd_DQ_in[51]\, \Sd_DQ_in[52]\, \Sd_DQ_in[53]\, 
        \Sd_DQ_in[54]\, \Sd_DQ_in[55]\, \Sd_DQ_in[56]\, 
        \Sd_DQ_in[57]\, \Sd_DQ_in[58]\, \Sd_DQ_in[59]\, 
        \Sd_DQ_in[60]\, \Sd_DQ_in[61]\, \Sd_DQ_in[62]\, 
        \Sd_DQ_in[63]\, \Sd_DQ_in[64]\, \Sd_DQ_in[65]\, 
        \Sd_DQ_in[66]\, \Sd_DQ_in[67]\, \Sd_DQ_in[68]\, 
        \Sd_DQ_in[69]\, \Sd_DQ_in[70]\, \Sd_DQ_in[71]\, 
        ExterCLk_c, CMOS_sample_c, mem_HL_c, Sync_X_c, Clock_Y_c, 
        spi_data_c, Clock_X_c, Sync_Y_c, spi_clock_c, Sh_co_c, 
        precharge_c, NoRowSel_c, CMOS_reset_c, Pre_co_c, 
        spi_load_c, SD_ras_n_c, SD_cas_n_c, SD_we_n_c, LVDS_O_c, 
        tok_c, DRY_c_c, \SD_cke_c_c[0]\, \SD_cs_n_c_c[1]\, 
        \SD_Clk_c_c[1]\, \SD_dqm_c_c_c_c_c_c_c_c[1]\, 
        \SD_addr_c[0]\, \SD_addr_c[1]\, \SD_addr_c[2]\, 
        \SD_addr_c[3]\, \SD_addr_c[4]\, \SD_addr_c[5]\, 
        \SD_addr_c[6]\, \SD_addr_c[7]\, \SD_addr_c[8]\, 
        \SD_addr_c[9]\, \SD_addr_c[10]\, \SD_addr_c[11]\, 
        \SD_addr_c[12]\, \GND\, \Counter_ref_0.refenlto5\, 
        \Main_ctl4SD_0.un6_sdramenreg\, CMOS_DrvX_0_AdcEn, 
        \intData2acc_RNIVOQA[0]\, \intData2acc_RNI2BV9[18]\, 
        \intData2acc_RNI6JV9[36]\, \intData2acc_RNIARV9[54]\, 
        \intData2acc_RNIBRV9[55]\, \intData2acc_RNI0TQA[1]\, 
        \intData2acc_RNI3BV9[19]\, \intData2acc_RNI7JV9[37]\, 
        \intData2acc_RNI11RA[2]\, \intData2acc_RNITEV9[20]\, 
        Sdram_ctl_v2_0_SD_rdEn_i, Sdram_ctl_v2_0_SD_wrEn_i, 
        FrameMk_0_LVDS_ok_i, Sdram_ini_0_Sd_iniOK_i, 
        \Sdram_cmd_0.N_264_0\, \Sdram_cmd_0.N_264_1\, 
        \Sdram_cmd_0.N_264_2\, CMOS_DrvX_0_SDramEn_0, 
        CMOS_DrvX_0_SDramEn_1, CMOS_DrvX_0_SDramEn_2, 
        CMOS_DrvX_0_SDramEn_3, CMOS_DrvX_0_SDramEn_4, 
        CMOS_DrvX_0_SDramEn_5, CMOS_DrvX_0_LVDSen_0, 
        CMOS_DrvX_0_LVDSen_1, CMOS_DrvX_0_LVDSen_2, 
        CMOS_DrvX_0_LVDSen_3, Main_ctl4SD_0_fifo_rst_n_0, 
        Main_ctl4SD_0_fifo_rst_n_1, Main_ctl4SD_0_fifo_rst_n_2, 
        Main_ctl4SD_0_fifo_rst_n_3, Main_ctl4SD_0_fifo_rst_n_4, 
        Main_ctl4SD_0_fifo_rst_n_5, Main_ctl4SD_0_fifo_rst_n_6, 
        GND_0, VCC_0 : std_logic;

    for all : FrameMk
	Use entity work.FrameMk(DEF_ARCH);
    for all : My_adder0_1
	Use entity work.My_adder0_1(DEF_ARCH);
    for all : Fifo_rd
	Use entity work.Fifo_rd(DEF_ARCH);
    for all : CMOS_DrvX
	Use entity work.CMOS_DrvX(DEF_ARCH);
    for all : My_adder0
	Use entity work.My_adder0(DEF_ARCH);
    for all : SDRAM_wr
	Use entity work.SDRAM_wr(DEF_ARCH);
    for all : Counter_ref
	Use entity work.Counter_ref(DEF_ARCH);
    for all : My_adder0_3
	Use entity work.My_adder0_3(DEF_ARCH);
    for all : SDRAM_Ref
	Use entity work.SDRAM_Ref(DEF_ARCH);
    for all : Sdram_cmd
	Use entity work.Sdram_cmd(DEF_ARCH);
    for all : Sdram_ini
	Use entity work.Sdram_ini(DEF_ARCH);
    for all : SDram_rd
	Use entity work.SDram_rd(DEF_ARCH);
    for all : Main_ctl4SD
	Use entity work.Main_ctl4SD(DEF_ARCH);
    for all : Fifo_rd_1
	Use entity work.Fifo_rd_1(DEF_ARCH);
    for all : Sdram_data
	Use entity work.Sdram_data(DEF_ARCH);
    for all : adc_muxtmp_test
	Use entity work.adc_muxtmp_test(DEF_ARCH);
    for all : PLL_Test1
	Use entity work.PLL_Test1(DEF_ARCH);
    for all : Sdram_ctl_v2
	Use entity work.Sdram_ctl_v2(DEF_ARCH);
    for all : My_adder0_2
	Use entity work.My_adder0_2(DEF_ARCH);
begin 


    \Sd_DQ_pad[28]\ : BIBUF
      port map(PAD => Sd_DQ(28), D => \Fifo_wr_0_Q_[28]\, E => 
        \Sdram_cmd_0.N_264_1\, Y => \Sd_DQ_in[28]\);
    
    \Sd_DQ_pad[62]\ : BIBUF
      port map(PAD => Sd_DQ(62), D => \Fifo_wr_0_Q_[62]\, E => 
        \Sdram_cmd_0.N_264\, Y => \Sd_DQ_in[62]\);
    
    \SD_cs_n_pad[1]\ : OUTBUF
      port map(D => \SD_cs_n_c_c[1]\, PAD => SD_cs_n(1));
    
    FrameMk_0 : FrameMk
      port map(FrameMk_GND => \GND\, CMOS_DrvX_0_LVDSen_3 => 
        CMOS_DrvX_0_LVDSen_3, FrameMk_VCC => \VCC\, 
        CMOS_DrvX_0_LVDSen => CMOS_DrvX_0_LVDSen, tok_c => tok_c, 
        LVDS_O_c => LVDS_O_c, Main_ctl4SD_0_ByteRdEn => 
        Main_ctl4SD_0_ByteRdEn, CMOS_DrvX_0_LVDSen_2 => 
        CMOS_DrvX_0_LVDSen_2, CMOS_DrvX_0_LVDSen_1 => 
        CMOS_DrvX_0_LVDSen_1, CMOS_DrvX_0_LVDSen_0 => 
        CMOS_DrvX_0_LVDSen_0, FrameMk_0_LVDS_ok => 
        FrameMk_0_LVDS_ok, FrameMk_0_LVDS_ok_i => 
        FrameMk_0_LVDS_ok_i, PLL_Test1_0_SysRst_O => 
        PLL_Test1_0_SysRst_O, PLL_Test1_0_Sys_66M_Clk => 
        PLL_Test1_0_Sys_66M_Clk);
    
    Sync_Y_pad : OUTBUF
      port map(D => Sync_Y_c, PAD => Sync_Y);
    
    \Sd_DQ_pad[47]\ : BIBUF
      port map(PAD => Sd_DQ(47), D => \Fifo_wr_0_Q_[47]\, E => 
        \Sdram_cmd_0.N_264_2\, Y => \Sd_DQ_in[47]\);
    
    \SD_ba_pad[0]\ : OUTBUF
      port map(D => \GND\, PAD => SD_ba(0));
    
    \My_adder0_3\ : My_adder0_1
      port map(intData2acc_RNIEVV9(64) => 
        \intData2acc_RNIEVV9[64]\, intData2acc_RNIDVV9(63) => 
        \intData2acc_RNIDVV9[63]\, intData2acc_RNIGVV9(66) => 
        \intData2acc_RNIGVV9[66]\, intData2acc_RNIDRV9(56) => 
        \intData2acc_RNIDRV9[56]\, intData2acc_RNIERV9(57) => 
        \intData2acc_RNIERV9[57]\, intData2acc_RNIHVV9(67) => 
        \intData2acc_RNIHVV9[67]\, intData2acc_RNIAVV9(60) => 
        \intData2acc_RNIAVV9[60]\, intData2acc_RNIBVV9(61) => 
        \intData2acc_RNIBVV9[61]\, intData2acc_RNIFVV9(65) => 
        \intData2acc_RNIFVV9[65]\, intData2acc_RNIPB46(71) => 
        \intData2acc_RNIPB46[71]\, intData2acc_RNIGRV9(59) => 
        \intData2acc_RNIGRV9[59]\, intData2acc_RNIGRV9(58) => 
        \intData2acc_RNIGRV9[58]\, intData2acc_RNICVV9(62) => 
        \intData2acc_RNICVV9[62]\, intData2acc_RNID30A(70) => 
        \intData2acc_RNID30A[70]\, intData2acc_RNIARV9(54) => 
        \intData2acc_RNIARV9[54]\, intData2acc_RNIBRV9(55) => 
        \intData2acc_RNIBRV9[55]\, \Z\\My_adder0_3_Sum_[15]\\\
         => \My_adder0_3_Sum_[15]\, \Z\\My_adder0_3_Sum_[12]\\\
         => \My_adder0_3_Sum_[12]\, \Z\\My_adder0_3_Sum_[6]\\\
         => \My_adder0_3_Sum_[6]\, \Z\\My_adder0_3_Sum_[10]\\\
         => \My_adder0_3_Sum_[10]\, \Z\\My_adder0_3_Sum_[9]\\\
         => \My_adder0_3_Sum_[9]\, \Z\\My_adder0_3_Sum_[7]\\\ => 
        \My_adder0_3_Sum_[7]\, N_6 => \Main_ctl4SD_0.N_6\, 
        \Z\\My_adder0_3_Sum_[11]\\\ => \My_adder0_3_Sum_[11]\, 
        \Z\\My_adder0_3_Sum_[1]\\\ => \My_adder0_3_Sum_[1]\, 
        \Z\\My_adder0_3_Sum_[3]\\\ => \My_adder0_3_Sum_[3]\, 
        \Z\\My_adder0_3_Sum_[13]\\\ => \My_adder0_3_Sum_[13]\, 
        \Z\\My_adder0_3_Sum_[0]\\\ => \My_adder0_3_Sum_[0]\, 
        \Z\\My_adder0_3_Sum_[8]\\\ => \My_adder0_3_Sum_[8]\, 
        \Z\\My_adder0_3_Sum_[14]\\\ => \My_adder0_3_Sum_[14]\, 
        \Z\\My_adder0_3_Sum_[2]\\\ => \My_adder0_3_Sum_[2]\, 
        \Z\\My_adder0_3_Sum_[4]\\\ => \My_adder0_3_Sum_[4]\, N_4
         => \Main_ctl4SD_0.N_4\, \Z\\My_adder0_3_Sum_[5]\\\ => 
        \My_adder0_3_Sum_[5]\, \Z\\My_adder0_3_Sum_[17]\\\ => 
        \My_adder0_3_Sum_[17]\, My_adder0_1_GND => \GND\, 
        \Z\\My_adder0_3_Sum_[16]\\\ => \My_adder0_3_Sum_[16]\, 
        \Z\\adc_muxtmp_test_0_DataOut55to42_[43]\\\ => 
        \adc_muxtmp_test_0_DataOut55to42_[43]\);
    
    \Sd_DQ_pad[69]\ : BIBUF
      port map(PAD => Sd_DQ(69), D => \Fifo_wr_0_Q_[69]\, E => 
        \Sdram_cmd_0.N_264\, Y => \Sd_DQ_in[69]\);
    
    \Sd_DQ_pad[66]\ : BIBUF
      port map(PAD => Sd_DQ(66), D => \Fifo_wr_0_Q_[66]\, E => 
        \Sdram_cmd_0.N_264\, Y => \Sd_DQ_in[66]\);
    
    \Sd_DQ_pad[32]\ : BIBUF
      port map(PAD => Sd_DQ(32), D => \Fifo_wr_0_Q_[32]\, E => 
        \Sdram_cmd_0.N_264_1\, Y => \Sd_DQ_in[32]\);
    
    Fifo_wr_0 : Fifo_rd
      port map(\Z\\Fifo_wr_0_Q_[27]\\\ => \Fifo_wr_0_Q_[27]\, 
        \Z\\Fifo_wr_0_Q_[23]\\\ => \Fifo_wr_0_Q_[23]\, 
        \Z\\Fifo_wr_0_Q_[69]\\\ => \Fifo_wr_0_Q_[69]\, 
        \Z\\Fifo_wr_0_Q_[1]\\\ => \Fifo_wr_0_Q_[1]\, 
        \Z\\Fifo_wr_0_Q_[67]\\\ => \Fifo_wr_0_Q_[67]\, 
        \Z\\Fifo_wr_0_Q_[4]\\\ => \Fifo_wr_0_Q_[4]\, 
        \Z\\Fifo_wr_0_Q_[63]\\\ => \Fifo_wr_0_Q_[63]\, 
        \Z\\Fifo_wr_0_Q_[7]\\\ => \Fifo_wr_0_Q_[7]\, 
        \Z\\Fifo_wr_0_Q_[56]\\\ => \Fifo_wr_0_Q_[56]\, 
        \Z\\Fifo_wr_0_Q_[25]\\\ => \Fifo_wr_0_Q_[25]\, 
        \Z\\Fifo_wr_0_Q_[24]\\\ => \Fifo_wr_0_Q_[24]\, 
        \Z\\Fifo_wr_0_Q_[48]\\\ => \Fifo_wr_0_Q_[48]\, 
        \Z\\Fifo_wr_0_Q_[65]\\\ => \Fifo_wr_0_Q_[65]\, 
        \Z\\Fifo_wr_0_Q_[64]\\\ => \Fifo_wr_0_Q_[64]\, 
        \Z\\Fifo_wr_0_Q_[51]\\\ => \Fifo_wr_0_Q_[51]\, 
        \Z\\Fifo_wr_0_Q_[38]\\\ => \Fifo_wr_0_Q_[38]\, 
        \Z\\Fifo_wr_0_Q_[71]\\\ => \Fifo_wr_0_Q_[71]\, 
        \Z\\Fifo_wr_0_Q_[50]\\\ => \Fifo_wr_0_Q_[50]\, 
        \Z\\Fifo_wr_0_Q_[70]\\\ => \Fifo_wr_0_Q_[70]\, 
        \Z\\Fifo_wr_0_Q_[18]\\\ => \Fifo_wr_0_Q_[18]\, 
        \Z\\Fifo_wr_0_Q_[6]\\\ => \Fifo_wr_0_Q_[6]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[71]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[71]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[70]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[70]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[69]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[69]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[68]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[68]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[67]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[67]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[66]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[66]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[65]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[65]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[64]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[64]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[63]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[63]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[62]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[62]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[61]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[61]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[60]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[60]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[59]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[59]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[58]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[58]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[57]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[57]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[56]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[56]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[55]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[55]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[54]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[54]\, \Z\\Fifo_wr_0_Q_[46]\\\
         => \Fifo_wr_0_Q_[46]\, \Z\\Fifo_wr_0_Q_[52]\\\ => 
        \Fifo_wr_0_Q_[52]\, \Z\\Fifo_wr_0_Q_[36]\\\ => 
        \Fifo_wr_0_Q_[36]\, \Z\\Fifo_wr_0_Q_[59]\\\ => 
        \Fifo_wr_0_Q_[59]\, \Z\\Fifo_wr_0_Q_[0]\\\ => 
        \Fifo_wr_0_Q_[0]\, \Z\\Fifo_wr_0_Q_[16]\\\ => 
        \Fifo_wr_0_Q_[16]\, \Z\\Fifo_wr_0_Q_[57]\\\ => 
        \Fifo_wr_0_Q_[57]\, \Z\\Fifo_wr_0_Q_[41]\\\ => 
        \Fifo_wr_0_Q_[41]\, \Z\\Fifo_wr_0_Q_[53]\\\ => 
        \Fifo_wr_0_Q_[53]\, \Z\\Fifo_wr_0_Q_[40]\\\ => 
        \Fifo_wr_0_Q_[40]\, Sdram_cmd_0_WFifo_re => 
        Sdram_cmd_0_WFifo_re, \Z\\Fifo_wr_0_Q_[31]\\\ => 
        \Fifo_wr_0_Q_[31]\, \Z\\Fifo_wr_0_Q_[28]\\\ => 
        \Fifo_wr_0_Q_[28]\, \Z\\Fifo_wr_0_Q_[30]\\\ => 
        \Fifo_wr_0_Q_[30]\, \Z\\Fifo_wr_0_Q_[42]\\\ => 
        \Fifo_wr_0_Q_[42]\, \Z\\Fifo_wr_0_Q_[11]\\\ => 
        \Fifo_wr_0_Q_[11]\, \Z\\Fifo_wr_0_Q_[10]\\\ => 
        \Fifo_wr_0_Q_[10]\, \Z\\Fifo_wr_0_Q_[55]\\\ => 
        \Fifo_wr_0_Q_[55]\, \Z\\Fifo_wr_0_Q_[68]\\\ => 
        \Fifo_wr_0_Q_[68]\, \Z\\Fifo_wr_0_Q_[54]\\\ => 
        \Fifo_wr_0_Q_[54]\, \Z\\Fifo_wr_0_Q_[49]\\\ => 
        \Fifo_wr_0_Q_[49]\, \Z\\Fifo_wr_0_Q_[9]\\\ => 
        \Fifo_wr_0_Q_[9]\, \Z\\Fifo_wr_0_Q_[5]\\\ => 
        \Fifo_wr_0_Q_[5]\, Fifo_wr_0_AFULL => Fifo_wr_0_AFULL, 
        \Z\\Fifo_wr_0_Q_[32]\\\ => \Fifo_wr_0_Q_[32]\, 
        \Z\\Fifo_wr_0_Q_[47]\\\ => \Fifo_wr_0_Q_[47]\, 
        \Z\\Fifo_wr_0_Q_[43]\\\ => \Fifo_wr_0_Q_[43]\, 
        Main_ctl4SD_0_fifo_rst_n_3 => Main_ctl4SD_0_fifo_rst_n_3, 
        \Z\\Fifo_wr_0_Q_[12]\\\ => \Fifo_wr_0_Q_[12]\, 
        Main_ctl4SD_0_Fifo_wr => Main_ctl4SD_0_Fifo_wr, 
        \Z\\Fifo_wr_0_Q_[26]\\\ => \Fifo_wr_0_Q_[26]\, 
        \Z\\Fifo_wr_0_Q_[39]\\\ => \Fifo_wr_0_Q_[39]\, 
        \Z\\Fifo_wr_0_Q_[19]\\\ => \Fifo_wr_0_Q_[19]\, 
        \Z\\Fifo_wr_0_Q_[37]\\\ => \Fifo_wr_0_Q_[37]\, 
        \Z\\Fifo_wr_0_Q_[3]\\\ => \Fifo_wr_0_Q_[3]\, 
        \Z\\Fifo_wr_0_Q_[33]\\\ => \Fifo_wr_0_Q_[33]\, 
        \Z\\Fifo_wr_0_Q_[66]\\\ => \Fifo_wr_0_Q_[66]\, 
        \Z\\Fifo_wr_0_Q_[17]\\\ => \Fifo_wr_0_Q_[17]\, 
        \Z\\Fifo_wr_0_Q_[13]\\\ => \Fifo_wr_0_Q_[13]\, 
        \Z\\Fifo_wr_0_Q_[45]\\\ => \Fifo_wr_0_Q_[45]\, 
        \Z\\Fifo_wr_0_Q_[44]\\\ => \Fifo_wr_0_Q_[44]\, 
        \Z\\Fifo_wr_0_Q_[21]\\\ => \Fifo_wr_0_Q_[21]\, 
        \Z\\Fifo_wr_0_Q_[2]\\\ => \Fifo_wr_0_Q_[2]\, 
        \Z\\Fifo_wr_0_Q_[20]\\\ => \Fifo_wr_0_Q_[20]\, 
        \Z\\Fifo_wr_0_Q_[61]\\\ => \Fifo_wr_0_Q_[61]\, 
        \Z\\Fifo_wr_0_Q_[35]\\\ => \Fifo_wr_0_Q_[35]\, 
        \Z\\Fifo_wr_0_Q_[34]\\\ => \Fifo_wr_0_Q_[34]\, 
        \Z\\Fifo_wr_0_Q_[60]\\\ => \Fifo_wr_0_Q_[60]\, 
        \Z\\Fifo_wr_0_Q_[15]\\\ => \Fifo_wr_0_Q_[15]\, 
        \Z\\Fifo_wr_0_Q_[14]\\\ => \Fifo_wr_0_Q_[14]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[35]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[35]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[34]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[34]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[33]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[33]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[32]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[32]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[31]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[31]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[30]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[30]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[29]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[29]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[28]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[28]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[27]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[27]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[26]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[26]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[25]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[25]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[24]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[24]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[23]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[23]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[22]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[22]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[21]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[21]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[20]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[20]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[19]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[19]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[18]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[18]\, 
        Main_ctl4SD_0_fifo_rst_n_4 => Main_ctl4SD_0_fifo_rst_n_4, 
        \Z\\Fifo_wr_0_Q_[22]\\\ => \Fifo_wr_0_Q_[22]\, 
        \Z\\Fifo_wr_0_Q_[8]\\\ => \Fifo_wr_0_Q_[8]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[53]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[53]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[52]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[52]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[51]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[51]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[50]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[50]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[49]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[49]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[48]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[48]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[47]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[47]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[46]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[46]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[45]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[45]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[44]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[44]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[43]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[43]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[42]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[42]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[41]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[41]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[40]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[40]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[39]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[39]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[38]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[38]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[37]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[37]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[36]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[36]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[17]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[17]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[16]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[16]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[15]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[15]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[14]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[14]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[13]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[13]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[12]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[12]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[11]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[11]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[10]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[10]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[9]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[9]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[8]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[8]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[7]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[7]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[6]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[6]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[5]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[5]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[4]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[4]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[3]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[3]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[2]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[2]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[1]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[1]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[0]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[0]\, Fifo_rd_VCC => \VCC\, 
        Main_ctl4SD_0_fifo_rst_n => Main_ctl4SD_0_fifo_rst_n, 
        \Z\\Fifo_wr_0_Q_[62]\\\ => \Fifo_wr_0_Q_[62]\, 
        Main_ctl4SD_0_fifo_rst_n_5 => Main_ctl4SD_0_fifo_rst_n_5, 
        \Z\\Fifo_wr_0_Q_[29]\\\ => \Fifo_wr_0_Q_[29]\, 
        Main_ctl4SD_0_fifo_rst_n_6 => Main_ctl4SD_0_fifo_rst_n_6, 
        PLL_Test1_0_Sys_66M_Clk => PLL_Test1_0_Sys_66M_Clk, 
        \Z\\Fifo_wr_0_Q_[58]\\\ => \Fifo_wr_0_Q_[58]\, 
        Fifo_rd_GND => \GND\);
    
    \Sd_DQ_pad[11]\ : BIBUF
      port map(PAD => Sd_DQ(11), D => \Fifo_wr_0_Q_[11]\, E => 
        \Sdram_cmd_0.N_264_0\, Y => \Sd_DQ_in[11]\);
    
    SD_cas_n_pad : OUTBUF
      port map(D => SD_cas_n_c, PAD => SD_cas_n);
    
    CMOS_reset_pad : OUTBUF
      port map(D => CMOS_reset_c, PAD => CMOS_reset);
    
    \Sd_DQ_pad[60]\ : BIBUF
      port map(PAD => Sd_DQ(60), D => \Fifo_wr_0_Q_[60]\, E => 
        \Sdram_cmd_0.N_264\, Y => \Sd_DQ_in[60]\);
    
    Sh_co_pad : OUTBUF
      port map(D => Sh_co_c, PAD => Sh_co);
    
    \Sd_DQ_pad[21]\ : BIBUF
      port map(PAD => Sd_DQ(21), D => \Fifo_wr_0_Q_[21]\, E => 
        \Sdram_cmd_0.N_264_0\, Y => \Sd_DQ_in[21]\);
    
    \Sd_DQ_pad[39]\ : BIBUF
      port map(PAD => Sd_DQ(39), D => \Fifo_wr_0_Q_[39]\, E => 
        \Sdram_cmd_0.N_264_1\, Y => \Sd_DQ_in[39]\);
    
    \Sd_DQ_pad[36]\ : BIBUF
      port map(PAD => Sd_DQ(36), D => \Fifo_wr_0_Q_[36]\, E => 
        \Sdram_cmd_0.N_264_1\, Y => \Sd_DQ_in[36]\);
    
    \Sd_DQ_pad[2]\ : BIBUF
      port map(PAD => Sd_DQ(2), D => \Fifo_wr_0_Q_[2]\, E => 
        \Sdram_cmd_0.N_264_1\, Y => \Sd_DQ_in[2]\);
    
    CMOS_DrvX_0 : CMOS_DrvX
      port map(CMOS_reset_c => CMOS_reset_c, CMOS_sample_c => 
        CMOS_sample_c, precharge_c => precharge_c, mem_HL_c => 
        mem_HL_c, spi_load_c => spi_load_c, spi_data_c => 
        spi_data_c, spi_clock_c => spi_clock_c, CMOS_DrvX_VCC => 
        \VCC\, PLL_Test1_0_ADC_66M_Clk => PLL_Test1_0_ADC_66M_Clk, 
        DRY_c_c => DRY_c_c, CMOS_DrvX_0_AdcEn => 
        CMOS_DrvX_0_AdcEn, Sync_Y_c => Sync_Y_c, Clock_Y_c => 
        Clock_Y_c, NoRowSel_c => NoRowSel_c, Pre_co_c => Pre_co_c, 
        Sh_co_c => Sh_co_c, Sync_X_c => Sync_X_c, Clock_X_c => 
        Clock_X_c, CMOS_DrvX_0_LVDSen_3 => CMOS_DrvX_0_LVDSen_3, 
        PLL_Test1_0_Sys_66M_Clk => PLL_Test1_0_Sys_66M_Clk, 
        PLL_Test1_0_SysRst_O => PLL_Test1_0_SysRst_O, 
        CMOS_DrvX_0_LVDSen_2 => CMOS_DrvX_0_LVDSen_2, 
        CMOS_DrvX_0_LVDSen_1 => CMOS_DrvX_0_LVDSen_1, 
        CMOS_DrvX_0_LVDSen_0 => CMOS_DrvX_0_LVDSen_0, 
        CMOS_DrvX_0_SDramEn_5 => CMOS_DrvX_0_SDramEn_5, 
        CMOS_DrvX_0_SDramEn_4 => CMOS_DrvX_0_SDramEn_4, 
        CMOS_DrvX_0_SDramEn_3 => CMOS_DrvX_0_SDramEn_3, 
        CMOS_DrvX_0_SDramEn_2 => CMOS_DrvX_0_SDramEn_2, 
        CMOS_DrvX_0_SDramEn_1 => CMOS_DrvX_0_SDramEn_1, 
        CMOS_DrvX_0_SDramEn_0 => CMOS_DrvX_0_SDramEn_0, 
        Sdram_cmd_0_SDoneFrameOk => Sdram_cmd_0_SDoneFrameOk, 
        FrameMk_0_LVDS_ok => FrameMk_0_LVDS_ok, 
        CMOS_DrvX_0_LVDSen => CMOS_DrvX_0_LVDSen, 
        CMOS_DrvX_0_SDramEn => CMOS_DrvX_0_SDramEn, CMOS_DrvX_GND
         => \GND\);
    
    \SD_addr_pad[7]\ : OUTBUF
      port map(D => \SD_addr_c[7]\, PAD => SD_addr(7));
    
    \Sd_DQ_pad[30]\ : BIBUF
      port map(PAD => Sd_DQ(30), D => \Fifo_wr_0_Q_[30]\, E => 
        \Sdram_cmd_0.N_264_1\, Y => \Sd_DQ_in[30]\);
    
    \SD_cke_pad[1]\ : OUTBUF
      port map(D => \SD_cke_c_c[0]\, PAD => SD_cke(1));
    
    precharge_pad : OUTBUF
      port map(D => precharge_c, PAD => precharge);
    
    \My_adder0_2\ : My_adder0
      port map(intData2acc_RNICNV9(46) => 
        \intData2acc_RNICNV9[46]\, intData2acc_RNIBNV9(45) => 
        \intData2acc_RNIBNV9[45]\, intData2acc_RNI9RV9(51) => 
        \intData2acc_RNI9RV9[51]\, intData2acc_RNI6JV9(36) => 
        \intData2acc_RNI6JV9[36]\, intData2acc_RNI7JV9(37) => 
        \intData2acc_RNI7JV9[37]\, intData2acc_RNI6NV9(40) => 
        \intData2acc_RNI6NV9[40]\, intData2acc_RNIENV9(48) => 
        \intData2acc_RNIENV9[48]\, intData2acc_RNI8RV9(50) => 
        \intData2acc_RNI8RV9[50]\, intData2acc_RNIBJV9(38) => 
        \intData2acc_RNIBJV9[38]\, intData2acc_RNICJV9(39) => 
        \intData2acc_RNICJV9[39]\, intData2acc_RNIFNV9(49) => 
        \intData2acc_RNIFNV9[49]\, intData2acc_RNI8NV9(42) => 
        \intData2acc_RNI8NV9[42]\, intData2acc_RNI9NV9(43) => 
        \intData2acc_RNI9NV9[43]\, intData2acc_RNIDNV9(47) => 
        \intData2acc_RNIDNV9[47]\, intData2acc_RNI7NV9(41) => 
        \intData2acc_RNI7NV9[41]\, intData2acc_RNIANV9(44) => 
        \intData2acc_RNIANV9[44]\, intData2acc_RNIBRV9(53) => 
        \intData2acc_RNIBRV9[53]\, intData2acc_RNIBRV9(52) => 
        \intData2acc_RNIBRV9[52]\, \Z\\My_adder0_2_Sum_[15]\\\
         => \My_adder0_2_Sum_[15]\, \Z\\My_adder0_2_Sum_[12]\\\
         => \My_adder0_2_Sum_[12]\, \Z\\My_adder0_2_Sum_[6]\\\
         => \My_adder0_2_Sum_[6]\, \Z\\My_adder0_2_Sum_[10]\\\
         => \My_adder0_2_Sum_[10]\, \Z\\My_adder0_2_Sum_[9]\\\
         => \My_adder0_2_Sum_[9]\, \Z\\My_adder0_2_Sum_[7]\\\ => 
        \My_adder0_2_Sum_[7]\, \Z\\My_adder0_2_Sum_[11]\\\ => 
        \My_adder0_2_Sum_[11]\, \Z\\My_adder0_2_Sum_[1]\\\ => 
        \My_adder0_2_Sum_[1]\, \Z\\My_adder0_2_Sum_[3]\\\ => 
        \My_adder0_2_Sum_[3]\, \Z\\My_adder0_2_Sum_[13]\\\ => 
        \My_adder0_2_Sum_[13]\, \Z\\My_adder0_2_Sum_[0]\\\ => 
        \My_adder0_2_Sum_[0]\, \Z\\My_adder0_2_Sum_[8]\\\ => 
        \My_adder0_2_Sum_[8]\, \Z\\My_adder0_2_Sum_[14]\\\ => 
        \My_adder0_2_Sum_[14]\, 
        \Z\\adc_muxtmp_test_0_DataOut41to28_[29]\\\ => 
        \adc_muxtmp_test_0_DataOut41to28_[29]\, 
        \Z\\My_adder0_2_Sum_[2]\\\ => \My_adder0_2_Sum_[2]\, 
        \Z\\My_adder0_2_Sum_[4]\\\ => \My_adder0_2_Sum_[4]\, 
        \Z\\My_adder0_2_Sum_[5]\\\ => \My_adder0_2_Sum_[5]\, 
        \Z\\My_adder0_2_Sum_[17]\\\ => \My_adder0_2_Sum_[17]\, 
        My_adder0_GND => \GND\, \Z\\My_adder0_2_Sum_[16]\\\ => 
        \My_adder0_2_Sum_[16]\);
    
    \Sd_DQ_pad[68]\ : BIBUF
      port map(PAD => Sd_DQ(68), D => \Fifo_wr_0_Q_[68]\, E => 
        \Sdram_cmd_0.N_264\, Y => \Sd_DQ_in[68]\);
    
    \Sd_DQ_pad[57]\ : BIBUF
      port map(PAD => Sd_DQ(57), D => \Fifo_wr_0_Q_[57]\, E => 
        \Sdram_cmd_0.N_264_2\, Y => \Sd_DQ_in[57]\);
    
    AdcClk_pad : OUTBUF
      port map(D => DRY_c_c, PAD => AdcClk);
    
    \SD_addr_pad[8]\ : OUTBUF
      port map(D => \SD_addr_c[8]\, PAD => SD_addr(8));
    
    NoRowSel_pad : OUTBUF
      port map(D => NoRowSel_c, PAD => NoRowSel);
    
    \Sd_DQ_pad[13]\ : BIBUF
      port map(PAD => Sd_DQ(13), D => \Fifo_wr_0_Q_[13]\, E => 
        \Sdram_cmd_0.N_264_0\, Y => \Sd_DQ_in[13]\);
    
    \Sd_DQ_pad[3]\ : BIBUF
      port map(PAD => Sd_DQ(3), D => \Fifo_wr_0_Q_[3]\, E => 
        \Sdram_cmd_0.N_264_1\, Y => \Sd_DQ_in[3]\);
    
    \SD_addr_pad[0]\ : OUTBUF
      port map(D => \SD_addr_c[0]\, PAD => SD_addr(0));
    
    \Sd_DQ_pad[42]\ : BIBUF
      port map(PAD => Sd_DQ(42), D => \Fifo_wr_0_Q_[42]\, E => 
        \Sdram_cmd_0.N_264_1\, Y => \Sd_DQ_in[42]\);
    
    \Sd_DQ_pad[23]\ : BIBUF
      port map(PAD => Sd_DQ(23), D => \Fifo_wr_0_Q_[23]\, E => 
        \Sdram_cmd_0.N_264_0\, Y => \Sd_DQ_in[23]\);
    
    SD_we_n_pad : OUTBUF
      port map(D => SD_we_n_c, PAD => SD_we_n);
    
    \Sd_DQ_pad[38]\ : BIBUF
      port map(PAD => Sd_DQ(38), D => \Fifo_wr_0_Q_[38]\, E => 
        \Sdram_cmd_0.N_264_1\, Y => \Sd_DQ_in[38]\);
    
    spi_clock_pad : OUTBUF
      port map(D => spi_clock_c, PAD => spi_clock);
    
    \Sd_DQ_pad[4]\ : BIBUF
      port map(PAD => Sd_DQ(4), D => \Fifo_wr_0_Q_[4]\, E => 
        \Sdram_cmd_0.N_264_2\, Y => \Sd_DQ_in[4]\);
    
    \SD_dqm_pad[2]\ : OUTBUF
      port map(D => \SD_dqm_c_c_c_c_c_c_c_c[1]\, PAD => SD_dqm(2));
    
    \Sd_DQ_pad[49]\ : BIBUF
      port map(PAD => Sd_DQ(49), D => \Fifo_wr_0_Q_[49]\, E => 
        \Sdram_cmd_0.N_264_2\, Y => \Sd_DQ_in[49]\);
    
    \Sd_DQ_pad[61]\ : BIBUF
      port map(PAD => Sd_DQ(61), D => \Fifo_wr_0_Q_[61]\, E => 
        \Sdram_cmd_0.N_264\, Y => \Sd_DQ_in[61]\);
    
    \Sd_DQ_pad[46]\ : BIBUF
      port map(PAD => Sd_DQ(46), D => \Fifo_wr_0_Q_[46]\, E => 
        \Sdram_cmd_0.N_264_2\, Y => \Sd_DQ_in[46]\);
    
    GND_i : GND
      port map(Y => \GND\);
    
    \SD_addr_pad[4]\ : OUTBUF
      port map(D => \SD_addr_c[4]\, PAD => SD_addr(4));
    
    VCC_i_0 : VCC
      port map(Y => VCC_0);
    
    ExterCLk_pad : INBUF
      port map(PAD => ExterCLk, Y => ExterCLk_c);
    
    \Sd_DQ_pad[5]\ : BIBUF
      port map(PAD => Sd_DQ(5), D => \Fifo_wr_0_Q_[5]\, E => 
        \Sdram_cmd_0.N_264_2\, Y => \Sd_DQ_in[5]\);
    
    \Sd_DQ_pad[40]\ : BIBUF
      port map(PAD => Sd_DQ(40), D => \Fifo_wr_0_Q_[40]\, E => 
        \Sdram_cmd_0.N_264_1\, Y => \Sd_DQ_in[40]\);
    
    \SD_cs_n_pad[0]\ : OUTBUF
      port map(D => \SD_cs_n_c_c[1]\, PAD => SD_cs_n(0));
    
    Clock_X_pad : OUTBUF
      port map(D => Clock_X_c, PAD => Clock_X);
    
    \Sd_DQ_pad[31]\ : BIBUF
      port map(PAD => Sd_DQ(31), D => \Fifo_wr_0_Q_[31]\, E => 
        \Sdram_cmd_0.N_264_1\, Y => \Sd_DQ_in[31]\);
    
    \Sd_DQ_pad[15]\ : BIBUF
      port map(PAD => Sd_DQ(15), D => \Fifo_wr_0_Q_[15]\, E => 
        \Sdram_cmd_0.N_264_0\, Y => \Sd_DQ_in[15]\);
    
    \SD_addr_pad[2]\ : OUTBUF
      port map(D => \SD_addr_c[2]\, PAD => SD_addr(2));
    
    SDRAM_wr_0 : SDRAM_wr
      port map(\Z\\SDRAM_wr_0_wr_state_[2]\\\ => 
        \SDRAM_wr_0_wr_state_[2]\, \Z\\SDRAM_wr_0_wr_state_[1]\\\
         => \SDRAM_wr_0_wr_state_[1]\, 
        \Z\\SDRAM_wr_0_wr_state_[0]\\\ => 
        \SDRAM_wr_0_wr_state_[0]\, Sdram_ctl_v2_0_SD_wrEn_i => 
        Sdram_ctl_v2_0_SD_wrEn_i, PLL_Test1_0_SysRst_O => 
        PLL_Test1_0_SysRst_O, PLL_Test1_0_Sys_66M_Clk => 
        PLL_Test1_0_Sys_66M_Clk, SDRAM_wr_0_SD_WrOK => 
        SDRAM_wr_0_SD_WrOK, Sdram_cmd_0_wrrow_end => 
        Sdram_cmd_0_wrrow_end, Sdram_ctl_v2_0_SD_wrEn => 
        Sdram_ctl_v2_0_SD_wrEn);
    
    \Sd_DQ_pad[70]\ : BIBUF
      port map(PAD => Sd_DQ(70), D => \Fifo_wr_0_Q_[70]\, E => 
        \Sdram_cmd_0.N_264\, Y => \Sd_DQ_in[70]\);
    
    \Sd_DQ_pad[25]\ : BIBUF
      port map(PAD => Sd_DQ(25), D => \Fifo_wr_0_Q_[25]\, E => 
        \Sdram_cmd_0.N_264_0\, Y => \Sd_DQ_in[25]\);
    
    SD_ras_n_pad : OUTBUF
      port map(D => SD_ras_n_c, PAD => SD_ras_n);
    
    \Sd_DQ_pad[52]\ : BIBUF
      port map(PAD => Sd_DQ(52), D => \Fifo_wr_0_Q_[52]\, E => 
        \Sdram_cmd_0.N_264_2\, Y => \Sd_DQ_in[52]\);
    
    \Sd_DQ_pad[48]\ : BIBUF
      port map(PAD => Sd_DQ(48), D => \Fifo_wr_0_Q_[48]\, E => 
        \Sdram_cmd_0.N_264_2\, Y => \Sd_DQ_in[48]\);
    
    \Sd_DQ_pad[63]\ : BIBUF
      port map(PAD => Sd_DQ(63), D => \Fifo_wr_0_Q_[63]\, E => 
        \Sdram_cmd_0.N_264\, Y => \Sd_DQ_in[63]\);
    
    \Sd_DQ_pad[59]\ : BIBUF
      port map(PAD => Sd_DQ(59), D => \Fifo_wr_0_Q_[59]\, E => 
        \Sdram_cmd_0.N_264_2\, Y => \Sd_DQ_in[59]\);
    
    VCC_i : VCC
      port map(Y => \VCC\);
    
    \Sd_DQ_pad[14]\ : BIBUF
      port map(PAD => Sd_DQ(14), D => \Fifo_wr_0_Q_[14]\, E => 
        \Sdram_cmd_0.N_264_0\, Y => \Sd_DQ_in[14]\);
    
    \Sd_DQ_pad[56]\ : BIBUF
      port map(PAD => Sd_DQ(56), D => \Fifo_wr_0_Q_[56]\, E => 
        \Sdram_cmd_0.N_264_2\, Y => \Sd_DQ_in[56]\);
    
    Counter_ref_0 : Counter_ref
      port map(refenlto5 => \Counter_ref_0.refenlto5\, 
        Sdram_ctl_v2_0_SD_RefEn => Sdram_ctl_v2_0_SD_RefEn, 
        PLL_Test1_0_SysRst_O => PLL_Test1_0_SysRst_O, 
        PLL_Test1_0_Sys_66M_Clk => PLL_Test1_0_Sys_66M_Clk, 
        Main_ctl4SD_0_ByteRdEn => Main_ctl4SD_0_ByteRdEn, 
        CMOS_DrvX_0_LVDSen_2 => CMOS_DrvX_0_LVDSen_2);
    
    \Sd_DQ_pad[24]\ : BIBUF
      port map(PAD => Sd_DQ(24), D => \Fifo_wr_0_Q_[24]\, E => 
        \Sdram_cmd_0.N_264_0\, Y => \Sd_DQ_in[24]\);
    
    \SD_dqm_pad[4]\ : OUTBUF
      port map(D => \SD_dqm_c_c_c_c_c_c_c_c[1]\, PAD => SD_dqm(4));
    
    \Sd_DQ_pad[33]\ : BIBUF
      port map(PAD => Sd_DQ(33), D => \Fifo_wr_0_Q_[33]\, E => 
        \Sdram_cmd_0.N_264_1\, Y => \Sd_DQ_in[33]\);
    
    \SD_ba_pad[1]\ : OUTBUF
      port map(D => \GND\, PAD => SD_ba(1));
    
    \Sd_DQ_pad[50]\ : BIBUF
      port map(PAD => Sd_DQ(50), D => \Fifo_wr_0_Q_[50]\, E => 
        \Sdram_cmd_0.N_264_2\, Y => \Sd_DQ_in[50]\);
    
    \SD_Clk_pad[1]\ : OUTBUF
      port map(D => \SD_Clk_c_c[1]\, PAD => SD_Clk(1));
    
    \Sd_DQ_pad[41]\ : BIBUF
      port map(PAD => Sd_DQ(41), D => \Fifo_wr_0_Q_[41]\, E => 
        \Sdram_cmd_0.N_264_1\, Y => \Sd_DQ_in[41]\);
    
    My_adder0_0 : My_adder0_3
      port map(intData2acc_RNI6J36(10) => 
        \intData2acc_RNI6J36[10]\, intData2acc_RNIK507(9) => 
        \intData2acc_RNIK507[9]\, intData2acc_RNIBJ36(15) => 
        \intData2acc_RNIBJ36[15]\, intData2acc_RNIVOQA(0) => 
        \intData2acc_RNIVOQA[0]\, intData2acc_RNI0TQA(1) => 
        \intData2acc_RNI0TQA[1]\, intData2acc_RNIFHV6(4) => 
        \intData2acc_RNIFHV6[4]\, intData2acc_RNI8J36(12) => 
        \intData2acc_RNI8J36[12]\, intData2acc_RNIAJ36(14) => 
        \intData2acc_RNIAJ36[14]\, intData2acc_RNI11RA(2) => 
        \intData2acc_RNI11RA[2]\, intData2acc_RNIEDV6(3) => 
        \intData2acc_RNIEDV6[3]\, intData2acc_RNI9J36(13) => 
        \intData2acc_RNI9J36[13]\, intData2acc_RNIHPV6(6) => 
        \intData2acc_RNIHPV6[6]\, intData2acc_RNIITV6(7) => 
        \intData2acc_RNIITV6[7]\, intData2acc_RNI7J36(11) => 
        \intData2acc_RNI7J36[11]\, intData2acc_RNIDJ36(17) => 
        \intData2acc_RNIDJ36[17]\, intData2acc_RNIGLV6(5) => 
        \intData2acc_RNIGLV6[5]\, intData2acc_RNIJ107(8) => 
        \intData2acc_RNIJ107[8]\, intData2acc_RNICJ36(16) => 
        \intData2acc_RNICJ36[16]\, \Z\\My_adder0_0_Sum_[15]\\\
         => \My_adder0_0_Sum_[15]\, \Z\\My_adder0_0_Sum_[12]\\\
         => \My_adder0_0_Sum_[12]\, \Z\\My_adder0_0_Sum_[6]\\\
         => \My_adder0_0_Sum_[6]\, \Z\\My_adder0_0_Sum_[10]\\\
         => \My_adder0_0_Sum_[10]\, \Z\\My_adder0_0_Sum_[9]\\\
         => \My_adder0_0_Sum_[9]\, \Z\\My_adder0_0_Sum_[7]\\\ => 
        \My_adder0_0_Sum_[7]\, \Z\\My_adder0_0_Sum_[11]\\\ => 
        \My_adder0_0_Sum_[11]\, \Z\\My_adder0_0_Sum_[1]\\\ => 
        \My_adder0_0_Sum_[1]\, \Z\\My_adder0_0_Sum_[3]\\\ => 
        \My_adder0_0_Sum_[3]\, \Z\\My_adder0_0_Sum_[13]\\\ => 
        \My_adder0_0_Sum_[13]\, \Z\\My_adder0_0_Sum_[0]\\\ => 
        \My_adder0_0_Sum_[0]\, \Z\\My_adder0_0_Sum_[8]\\\ => 
        \My_adder0_0_Sum_[8]\, \Z\\My_adder0_0_Sum_[14]\\\ => 
        \My_adder0_0_Sum_[14]\, \Z\\My_adder0_0_Sum_[2]\\\ => 
        \My_adder0_0_Sum_[2]\, \Z\\My_adder0_0_Sum_[4]\\\ => 
        \My_adder0_0_Sum_[4]\, \Z\\My_adder0_0_Sum_[5]\\\ => 
        \My_adder0_0_Sum_[5]\, \Z\\My_adder0_0_Sum_[17]\\\ => 
        \My_adder0_0_Sum_[17]\, My_adder0_3_GND => \GND\, 
        \Z\\My_adder0_0_Sum_[16]\\\ => \My_adder0_0_Sum_[16]\);
    
    \Sd_DQ_pad[65]\ : BIBUF
      port map(PAD => Sd_DQ(65), D => \Fifo_wr_0_Q_[65]\, E => 
        \Sdram_cmd_0.N_264\, Y => \Sd_DQ_in[65]\);
    
    \Sd_DQ_pad[71]\ : BIBUF
      port map(PAD => Sd_DQ(71), D => \Fifo_wr_0_Q_[71]\, E => 
        \Sdram_cmd_0.N_264\, Y => \Sd_DQ_in[71]\);
    
    DRY_pad : OUTBUF
      port map(D => DRY_c_c, PAD => DRY);
    
    CMOS_sample_pad : OUTBUF
      port map(D => CMOS_sample_c, PAD => CMOS_sample);
    
    \Sd_DQ_pad[58]\ : BIBUF
      port map(PAD => Sd_DQ(58), D => \Fifo_wr_0_Q_[58]\, E => 
        \Sdram_cmd_0.N_264_2\, Y => \Sd_DQ_in[58]\);
    
    SDRAM_Ref_0 : SDRAM_Ref
      port map(\Z\\SDRAM_Ref_0_Ref_state_[2]\\\ => 
        \SDRAM_Ref_0_Ref_state_[2]\, 
        \Z\\SDRAM_Ref_0_Ref_state_[1]\\\ => 
        \SDRAM_Ref_0_Ref_state_[1]\, 
        \Z\\SDRAM_Ref_0_Ref_state_[0]\\\ => 
        \SDRAM_Ref_0_Ref_state_[0]\, ref_ok_1 => 
        \SDRAM_Ref_0.ref_ok_1\, PLL_Test1_0_SysRst_O => 
        PLL_Test1_0_SysRst_O, PLL_Test1_0_Sys_66M_Clk => 
        PLL_Test1_0_Sys_66M_Clk, ref_ok_2 => 
        \SDRAM_Ref_0.ref_ok_2\, Sdram_ctl_v2_0_SD_RefEn => 
        Sdram_ctl_v2_0_SD_RefEn, Sdram_ini_0_Sd_iniOK => 
        Sdram_ini_0_Sd_iniOK, refenlto5 => 
        \Counter_ref_0.refenlto5\, Sdram_ctl_v2_0_SD_pdEN => 
        Sdram_ctl_v2_0_SD_pdEN);
    
    \SD_dqm_pad[1]\ : OUTBUF
      port map(D => \SD_dqm_c_c_c_c_c_c_c_c[1]\, PAD => SD_dqm(1));
    
    Sdram_cmd_0 : Sdram_cmd
      port map(SD_cs_n_c_c(1) => \SD_cs_n_c_c[1]\, 
        SD_dqm_c_c_c_c_c_c_c_c(1) => \SD_dqm_c_c_c_c_c_c_c_c[1]\, 
        SD_cke_c_c(0) => \SD_cke_c_c[0]\, SD_Clk_c_c(1) => 
        \SD_Clk_c_c[1]\, SD_addr_c(12) => \SD_addr_c[12]\, 
        SD_addr_c(11) => \SD_addr_c[11]\, SD_addr_c(10) => 
        \SD_addr_c[10]\, SD_addr_c(9) => \SD_addr_c[9]\, 
        SD_addr_c(8) => \SD_addr_c[8]\, SD_addr_c(7) => 
        \SD_addr_c[7]\, SD_addr_c(6) => \SD_addr_c[6]\, 
        SD_addr_c(5) => \SD_addr_c[5]\, SD_addr_c(4) => 
        \SD_addr_c[4]\, SD_addr_c(3) => \SD_addr_c[3]\, 
        SD_addr_c(2) => \SD_addr_c[2]\, SD_addr_c(1) => 
        \SD_addr_c[1]\, SD_addr_c(0) => \SD_addr_c[0]\, 
        Sdram_cmd_0_RFifo_we => Sdram_cmd_0_RFifo_we, 
        Sdram_cmd_0_rdrow_end => Sdram_cmd_0_rdrow_end, 
        Sdram_cmd_0_WFifo_re => Sdram_cmd_0_WFifo_re, 
        Sdram_cmd_0_wrrow_end => Sdram_cmd_0_wrrow_end, 
        SD_ras_n_c => SD_ras_n_c, SD_we_n_c => SD_we_n_c, 
        SD_cas_n_c => SD_cas_n_c, CMOS_DrvX_0_LVDSen => 
        CMOS_DrvX_0_LVDSen, Sdram_cmd_0_SDoneFrameOk => 
        Sdram_cmd_0_SDoneFrameOk, CMOS_DrvX_0_SDramEn => 
        CMOS_DrvX_0_SDramEn, PLL_Test1_0_SysRst_O => 
        PLL_Test1_0_SysRst_O, PLL_Test1_0_Sys_66M_Clk => 
        PLL_Test1_0_Sys_66M_Clk, LVDS_enReg => 
        \Sdram_cmd_0.LVDS_enReg\, CMOS_DrvX_0_LVDSen_2 => 
        CMOS_DrvX_0_LVDSen_2, \Z\\Sdram_ini_0_ini_state_[0]\\\
         => \Sdram_ini_0_ini_state_[0]\, un6_sdramenreg => 
        \Main_ctl4SD_0.un6_sdramenreg\, N_264 => 
        \Sdram_cmd_0.N_264\, \Z\\SDRAM_Ref_0_Ref_state_[0]\\\ => 
        \SDRAM_Ref_0_Ref_state_[0]\, 
        \Z\\SDRAM_Ref_0_Ref_state_[2]\\\ => 
        \SDRAM_Ref_0_Ref_state_[2]\, 
        \Z\\SDRAM_Ref_0_Ref_state_[1]\\\ => 
        \SDRAM_Ref_0_Ref_state_[1]\, PLL_Test1_0_Sdram_clk => 
        PLL_Test1_0_Sdram_clk, \Z\\SDram_rd_0_rd_state_[1]\\\ => 
        \SDram_rd_0_rd_state_[1]\, \Z\\SDram_rd_0_rd_state_[2]\\\
         => \SDram_rd_0_rd_state_[2]\, 
        \Z\\SDram_rd_0_rd_state_[0]\\\ => 
        \SDram_rd_0_rd_state_[0]\, 
        \Z\\Sdram_ini_0_ini_state_[2]\\\ => 
        \Sdram_ini_0_ini_state_[2]\, 
        \Z\\Sdram_ini_0_ini_state_[1]\\\ => 
        \Sdram_ini_0_ini_state_[1]\, N_264_0 => 
        \Sdram_cmd_0.N_264_0\, N_264_1 => \Sdram_cmd_0.N_264_1\, 
        \Z\\SDRAM_wr_0_wr_state_[1]\\\ => 
        \SDRAM_wr_0_wr_state_[1]\, \Z\\SDRAM_wr_0_wr_state_[0]\\\
         => \SDRAM_wr_0_wr_state_[0]\, 
        \Z\\SDRAM_wr_0_wr_state_[2]\\\ => 
        \SDRAM_wr_0_wr_state_[2]\, N_264_2 => 
        \Sdram_cmd_0.N_264_2\);
    
    Sync_X_pad : OUTBUF
      port map(D => Sync_X_c, PAD => Sync_X);
    
    \Sd_DQ_pad[35]\ : BIBUF
      port map(PAD => Sd_DQ(35), D => \Fifo_wr_0_Q_[35]\, E => 
        \Sdram_cmd_0.N_264_1\, Y => \Sd_DQ_in[35]\);
    
    \SD_dqm_pad[5]\ : OUTBUF
      port map(D => \SD_dqm_c_c_c_c_c_c_c_c[1]\, PAD => SD_dqm(5));
    
    Prebus1_pad : OUTBUF
      port map(D => \GND\, PAD => Prebus1);
    
    \Sd_DQ_pad[43]\ : BIBUF
      port map(PAD => Sd_DQ(43), D => \Fifo_wr_0_Q_[43]\, E => 
        \Sdram_cmd_0.N_264_2\, Y => \Sd_DQ_in[43]\);
    
    \SD_cke_pad[0]\ : OUTBUF
      port map(D => \SD_cke_c_c[0]\, PAD => SD_cke(0));
    
    \Sd_DQ_pad[64]\ : BIBUF
      port map(PAD => Sd_DQ(64), D => \Fifo_wr_0_Q_[64]\, E => 
        \Sdram_cmd_0.N_264\, Y => \Sd_DQ_in[64]\);
    
    LVDS_O_pad : OUTBUF
      port map(D => LVDS_O_c, PAD => LVDS_O);
    
    \Sd_DQ_pad[1]\ : BIBUF
      port map(PAD => Sd_DQ(1), D => \Fifo_wr_0_Q_[1]\, E => 
        \Sdram_cmd_0.N_264_0\, Y => \Sd_DQ_in[1]\);
    
    Sdram_ini_0 : Sdram_ini
      port map(\Z\\Sdram_ini_0_ini_state_[2]\\\ => 
        \Sdram_ini_0_ini_state_[2]\, 
        \Z\\Sdram_ini_0_ini_state_[1]\\\ => 
        \Sdram_ini_0_ini_state_[1]\, 
        \Z\\Sdram_ini_0_ini_state_[0]\\\ => 
        \Sdram_ini_0_ini_state_[0]\, PLL_Test1_0_SysRst_O => 
        PLL_Test1_0_SysRst_O, PLL_Test1_0_Sys_66M_Clk => 
        PLL_Test1_0_Sys_66M_Clk, Sdram_ctl_v2_0_SD_iniEn => 
        Sdram_ctl_v2_0_SD_iniEn, Sdram_ini_0_Sd_iniOK => 
        Sdram_ini_0_Sd_iniOK, Sdram_ini_0_Sd_iniOK_i => 
        Sdram_ini_0_Sd_iniOK_i);
    
    mem_HL_pad : OUTBUF
      port map(D => mem_HL_c, PAD => mem_HL);
    
    \SD_addr_pad[3]\ : OUTBUF
      port map(D => \SD_addr_c[3]\, PAD => SD_addr(3));
    
    SDram_rd_0 : SDram_rd
      port map(\Z\\SDram_rd_0_rd_state_[2]\\\ => 
        \SDram_rd_0_rd_state_[2]\, \Z\\SDram_rd_0_rd_state_[1]\\\
         => \SDram_rd_0_rd_state_[1]\, 
        \Z\\SDram_rd_0_rd_state_[0]\\\ => 
        \SDram_rd_0_rd_state_[0]\, Sdram_ctl_v2_0_SD_rdEn_i => 
        Sdram_ctl_v2_0_SD_rdEn_i, PLL_Test1_0_SysRst_O => 
        PLL_Test1_0_SysRst_O, PLL_Test1_0_Sys_66M_Clk => 
        PLL_Test1_0_Sys_66M_Clk, SDram_rd_0_SD_RdOK => 
        SDram_rd_0_SD_RdOK, Sdram_ctl_v2_0_SD_rdEn => 
        Sdram_ctl_v2_0_SD_rdEn, Sdram_cmd_0_rdrow_end => 
        Sdram_cmd_0_rdrow_end, Sdram_ctl_v2_0_SD_rdEN_noact => 
        Sdram_ctl_v2_0_SD_rdEN_noact);
    
    \Sd_DQ_pad[51]\ : BIBUF
      port map(PAD => Sd_DQ(51), D => \Fifo_wr_0_Q_[51]\, E => 
        \Sdram_cmd_0.N_264_2\, Y => \Sd_DQ_in[51]\);
    
    Main_ctl4SD_0 : Main_ctl4SD
      port map(intData2acc_RNIPB46(71) => 
        \intData2acc_RNIPB46[71]\, intData2acc_RNIFHV6(4) => 
        \intData2acc_RNIFHV6[4]\, intData2acc_RNIEDV6(3) => 
        \intData2acc_RNIEDV6[3]\, intData2acc_RNIITV6(7) => 
        \intData2acc_RNIITV6[7]\, intData2acc_RNIHPV6(6) => 
        \intData2acc_RNIHPV6[6]\, intData2acc_RNIGLV6(5) => 
        \intData2acc_RNIGLV6[5]\, intData2acc_RNI6J36(10) => 
        \intData2acc_RNI6J36[10]\, intData2acc_RNIK507(9) => 
        \intData2acc_RNIK507[9]\, intData2acc_RNIJ107(8) => 
        \intData2acc_RNIJ107[8]\, intData2acc_RNI9J36(13) => 
        \intData2acc_RNI9J36[13]\, intData2acc_RNI8J36(12) => 
        \intData2acc_RNI8J36[12]\, intData2acc_RNI7J36(11) => 
        \intData2acc_RNI7J36[11]\, intData2acc_RNICJ36(16) => 
        \intData2acc_RNICJ36[16]\, intData2acc_RNIBJ36(15) => 
        \intData2acc_RNIBJ36[15]\, intData2acc_RNIAJ36(14) => 
        \intData2acc_RNIAJ36[14]\, intData2acc_RNIDJ36(17) => 
        \intData2acc_RNIDJ36[17]\, intData2acc_RNIBN36(22) => 
        \intData2acc_RNIBN36[22]\, intData2acc_RNIAN36(21) => 
        \intData2acc_RNIAN36[21]\, intData2acc_RNIEN36(25) => 
        \intData2acc_RNIEN36[25]\, intData2acc_RNIDN36(24) => 
        \intData2acc_RNIDN36[24]\, intData2acc_RNITJS7(23) => 
        \intData2acc_RNITJS7[23]\, intData2acc_RNI2KS7(28) => 
        \intData2acc_RNI2KS7[28]\, intData2acc_RNI1KS7(27) => 
        \intData2acc_RNI1KS7[27]\, intData2acc_RNI0KS7(26) => 
        \intData2acc_RNI0KS7[26]\, intData2acc_RNI4JV9(31) => 
        \intData2acc_RNI4JV9[31]\, intData2acc_RNI3JV9(30) => 
        \intData2acc_RNI3JV9[30]\, intData2acc_RNI9FV9(29) => 
        \intData2acc_RNI9FV9[29]\, intData2acc_RNI5JV9(32) => 
        \intData2acc_RNI5JV9[32]\, intData2acc_RNI8JV9(35) => 
        \intData2acc_RNI8JV9[35]\, intData2acc_RNI6NV9(40) => 
        \intData2acc_RNI6NV9[40]\, intData2acc_RNICJV9(39) => 
        \intData2acc_RNICJV9[39]\, intData2acc_RNIBJV9(38) => 
        \intData2acc_RNIBJV9[38]\, intData2acc_RNI9NV9(43) => 
        \intData2acc_RNI9NV9[43]\, intData2acc_RNI8NV9(42) => 
        \intData2acc_RNI8NV9[42]\, intData2acc_RNI7NV9(41) => 
        \intData2acc_RNI7NV9[41]\, intData2acc_RNICNV9(46) => 
        \intData2acc_RNICNV9[46]\, intData2acc_RNIBNV9(45) => 
        \intData2acc_RNIBNV9[45]\, intData2acc_RNIANV9(44) => 
        \intData2acc_RNIANV9[44]\, intData2acc_RNIFNV9(49) => 
        \intData2acc_RNIFNV9[49]\, intData2acc_RNIENV9(48) => 
        \intData2acc_RNIENV9[48]\, intData2acc_RNIDNV9(47) => 
        \intData2acc_RNIDNV9[47]\, intData2acc_RNI9RV9(51) => 
        \intData2acc_RNI9RV9[51]\, intData2acc_RNI8RV9(50) => 
        \intData2acc_RNI8RV9[50]\, intData2acc_RNIERV9(57) => 
        \intData2acc_RNIERV9[57]\, intData2acc_RNIDRV9(56) => 
        \intData2acc_RNIDRV9[56]\, intData2acc_RNIBVV9(61) => 
        \intData2acc_RNIBVV9[61]\, intData2acc_RNIAVV9(60) => 
        \intData2acc_RNIAVV9[60]\, intData2acc_RNIGRV9(59) => 
        \intData2acc_RNIGRV9[59]\, intData2acc_RNIGRV9(58) => 
        \intData2acc_RNIGRV9[58]\, intData2acc_RNIEVV9(64) => 
        \intData2acc_RNIEVV9[64]\, intData2acc_RNIDVV9(63) => 
        \intData2acc_RNIDVV9[63]\, intData2acc_RNICVV9(62) => 
        \intData2acc_RNICVV9[62]\, intData2acc_RNIHVV9(67) => 
        \intData2acc_RNIHVV9[67]\, intData2acc_RNIGVV9(66) => 
        \intData2acc_RNIGVV9[66]\, intData2acc_RNIFVV9(65) => 
        \intData2acc_RNIFVV9[65]\, intData2acc_RNID30A(70) => 
        \intData2acc_RNID30A[70]\, intData2acc_RNIVOQA(0) => 
        \intData2acc_RNIVOQA[0]\, intData2acc_RNI2BV9(18) => 
        \intData2acc_RNI2BV9[18]\, intData2acc_RNI6JV9_0 => 
        \intData2acc_RNI6JV9[33]\, intData2acc_RNI6JV9_3 => 
        \intData2acc_RNI6JV9[36]\, intData2acc_RNI0TQA(1) => 
        \intData2acc_RNI0TQA[1]\, intData2acc_RNI3BV9(19) => 
        \intData2acc_RNI3BV9[19]\, intData2acc_RNI7JV9_0 => 
        \intData2acc_RNI7JV9[34]\, intData2acc_RNI7JV9_3 => 
        \intData2acc_RNI7JV9[37]\, intData2acc_RNI11RA(2) => 
        \intData2acc_RNI11RA[2]\, intData2acc_RNITEV9(20) => 
        \intData2acc_RNITEV9[20]\, pr_state_ns(8) => 
        \Sdram_ctl_v2_0.pr_state_ns[8]\, intData2acc_RNIARV9(54)
         => \intData2acc_RNIARV9[54]\, intData2acc_RNIBRV9_0 => 
        \intData2acc_RNIBRV9[52]\, intData2acc_RNIBRV9_1 => 
        \intData2acc_RNIBRV9[53]\, intData2acc_RNIBRV9_3 => 
        \intData2acc_RNIBRV9[55]\, Main_ctl4SD_0_ByteRdEn => 
        Main_ctl4SD_0_ByteRdEn, CMOS_DrvX_0_LVDSen_1 => 
        CMOS_DrvX_0_LVDSen_1, CMOS_DrvX_0_LVDSen_2 => 
        CMOS_DrvX_0_LVDSen_2, Main_ctl4SD_0_Fifo_wr => 
        Main_ctl4SD_0_Fifo_wr, Main_ctl4SD_0_fifo_rd => 
        Main_ctl4SD_0_fifo_rd, \Z\\Fifo_rd_0_Q_[71]\\\ => 
        \Fifo_rd_0_Q_[71]\, \Z\\Fifo_rd_0_Q_[70]\\\ => 
        \Fifo_rd_0_Q_[70]\, \Z\\Fifo_rd_0_Q_[69]\\\ => 
        \Fifo_rd_0_Q_[69]\, \Z\\Fifo_rd_0_Q_[68]\\\ => 
        \Fifo_rd_0_Q_[68]\, \Z\\Fifo_rd_0_Q_[67]\\\ => 
        \Fifo_rd_0_Q_[67]\, \Z\\Fifo_rd_0_Q_[66]\\\ => 
        \Fifo_rd_0_Q_[66]\, \Z\\Fifo_rd_0_Q_[65]\\\ => 
        \Fifo_rd_0_Q_[65]\, \Z\\Fifo_rd_0_Q_[64]\\\ => 
        \Fifo_rd_0_Q_[64]\, \Z\\Fifo_rd_0_Q_[63]\\\ => 
        \Fifo_rd_0_Q_[63]\, \Z\\Fifo_rd_0_Q_[62]\\\ => 
        \Fifo_rd_0_Q_[62]\, \Z\\Fifo_rd_0_Q_[61]\\\ => 
        \Fifo_rd_0_Q_[61]\, \Z\\Fifo_rd_0_Q_[60]\\\ => 
        \Fifo_rd_0_Q_[60]\, \Z\\Fifo_rd_0_Q_[59]\\\ => 
        \Fifo_rd_0_Q_[59]\, \Z\\Fifo_rd_0_Q_[58]\\\ => 
        \Fifo_rd_0_Q_[58]\, \Z\\Fifo_rd_0_Q_[57]\\\ => 
        \Fifo_rd_0_Q_[57]\, \Z\\Fifo_rd_0_Q_[56]\\\ => 
        \Fifo_rd_0_Q_[56]\, \Z\\Fifo_rd_0_Q_[55]\\\ => 
        \Fifo_rd_0_Q_[55]\, \Z\\Fifo_rd_0_Q_[54]\\\ => 
        \Fifo_rd_0_Q_[54]\, \Z\\Fifo_rd_0_Q_[53]\\\ => 
        \Fifo_rd_0_Q_[53]\, \Z\\Fifo_rd_0_Q_[52]\\\ => 
        \Fifo_rd_0_Q_[52]\, \Z\\Fifo_rd_0_Q_[51]\\\ => 
        \Fifo_rd_0_Q_[51]\, \Z\\Fifo_rd_0_Q_[50]\\\ => 
        \Fifo_rd_0_Q_[50]\, \Z\\Fifo_rd_0_Q_[49]\\\ => 
        \Fifo_rd_0_Q_[49]\, \Z\\Fifo_rd_0_Q_[48]\\\ => 
        \Fifo_rd_0_Q_[48]\, \Z\\Fifo_rd_0_Q_[47]\\\ => 
        \Fifo_rd_0_Q_[47]\, \Z\\Fifo_rd_0_Q_[46]\\\ => 
        \Fifo_rd_0_Q_[46]\, \Z\\Fifo_rd_0_Q_[45]\\\ => 
        \Fifo_rd_0_Q_[45]\, \Z\\Fifo_rd_0_Q_[44]\\\ => 
        \Fifo_rd_0_Q_[44]\, \Z\\Fifo_rd_0_Q_[43]\\\ => 
        \Fifo_rd_0_Q_[43]\, \Z\\Fifo_rd_0_Q_[42]\\\ => 
        \Fifo_rd_0_Q_[42]\, \Z\\Fifo_rd_0_Q_[41]\\\ => 
        \Fifo_rd_0_Q_[41]\, \Z\\Fifo_rd_0_Q_[40]\\\ => 
        \Fifo_rd_0_Q_[40]\, \Z\\Fifo_rd_0_Q_[39]\\\ => 
        \Fifo_rd_0_Q_[39]\, \Z\\Fifo_rd_0_Q_[38]\\\ => 
        \Fifo_rd_0_Q_[38]\, \Z\\Fifo_rd_0_Q_[37]\\\ => 
        \Fifo_rd_0_Q_[37]\, \Z\\Fifo_rd_0_Q_[36]\\\ => 
        \Fifo_rd_0_Q_[36]\, \Z\\Fifo_rd_0_Q_[35]\\\ => 
        \Fifo_rd_0_Q_[35]\, \Z\\Fifo_rd_0_Q_[34]\\\ => 
        \Fifo_rd_0_Q_[34]\, \Z\\Fifo_rd_0_Q_[33]\\\ => 
        \Fifo_rd_0_Q_[33]\, \Z\\Fifo_rd_0_Q_[32]\\\ => 
        \Fifo_rd_0_Q_[32]\, \Z\\Fifo_rd_0_Q_[31]\\\ => 
        \Fifo_rd_0_Q_[31]\, \Z\\Fifo_rd_0_Q_[30]\\\ => 
        \Fifo_rd_0_Q_[30]\, \Z\\Fifo_rd_0_Q_[29]\\\ => 
        \Fifo_rd_0_Q_[29]\, \Z\\Fifo_rd_0_Q_[28]\\\ => 
        \Fifo_rd_0_Q_[28]\, \Z\\Fifo_rd_0_Q_[27]\\\ => 
        \Fifo_rd_0_Q_[27]\, \Z\\Fifo_rd_0_Q_[26]\\\ => 
        \Fifo_rd_0_Q_[26]\, \Z\\Fifo_rd_0_Q_[25]\\\ => 
        \Fifo_rd_0_Q_[25]\, \Z\\Fifo_rd_0_Q_[24]\\\ => 
        \Fifo_rd_0_Q_[24]\, \Z\\Fifo_rd_0_Q_[23]\\\ => 
        \Fifo_rd_0_Q_[23]\, \Z\\Fifo_rd_0_Q_[22]\\\ => 
        \Fifo_rd_0_Q_[22]\, \Z\\Fifo_rd_0_Q_[21]\\\ => 
        \Fifo_rd_0_Q_[21]\, \Z\\Fifo_rd_0_Q_[20]\\\ => 
        \Fifo_rd_0_Q_[20]\, \Z\\Fifo_rd_0_Q_[19]\\\ => 
        \Fifo_rd_0_Q_[19]\, \Z\\Fifo_rd_0_Q_[18]\\\ => 
        \Fifo_rd_0_Q_[18]\, \Z\\Fifo_rd_0_Q_[17]\\\ => 
        \Fifo_rd_0_Q_[17]\, \Z\\Fifo_rd_0_Q_[16]\\\ => 
        \Fifo_rd_0_Q_[16]\, \Z\\Fifo_rd_0_Q_[15]\\\ => 
        \Fifo_rd_0_Q_[15]\, \Z\\Fifo_rd_0_Q_[14]\\\ => 
        \Fifo_rd_0_Q_[14]\, \Z\\Fifo_rd_0_Q_[13]\\\ => 
        \Fifo_rd_0_Q_[13]\, \Z\\Fifo_rd_0_Q_[12]\\\ => 
        \Fifo_rd_0_Q_[12]\, \Z\\Fifo_rd_0_Q_[11]\\\ => 
        \Fifo_rd_0_Q_[11]\, \Z\\Fifo_rd_0_Q_[10]\\\ => 
        \Fifo_rd_0_Q_[10]\, \Z\\Fifo_rd_0_Q_[9]\\\ => 
        \Fifo_rd_0_Q_[9]\, \Z\\Fifo_rd_0_Q_[8]\\\ => 
        \Fifo_rd_0_Q_[8]\, \Z\\Fifo_rd_0_Q_[7]\\\ => 
        \Fifo_rd_0_Q_[7]\, \Z\\Fifo_rd_0_Q_[6]\\\ => 
        \Fifo_rd_0_Q_[6]\, \Z\\Fifo_rd_0_Q_[5]\\\ => 
        \Fifo_rd_0_Q_[5]\, \Z\\Fifo_rd_0_Q_[4]\\\ => 
        \Fifo_rd_0_Q_[4]\, \Z\\Fifo_rd_0_Q_[3]\\\ => 
        \Fifo_rd_0_Q_[3]\, \Z\\Fifo_rd_0_Q_[2]\\\ => 
        \Fifo_rd_0_Q_[2]\, \Z\\Fifo_rd_0_Q_[1]\\\ => 
        \Fifo_rd_0_Q_[1]\, \Z\\Fifo_rd_0_Q_[0]\\\ => 
        \Fifo_rd_0_Q_[0]\, CMOS_DrvX_0_SDramEn_2 => 
        CMOS_DrvX_0_SDramEn_2, CMOS_DrvX_0_SDramEn_1 => 
        CMOS_DrvX_0_SDramEn_1, CMOS_DrvX_0_SDramEn => 
        CMOS_DrvX_0_SDramEn, CMOS_DrvX_0_SDramEn_5 => 
        CMOS_DrvX_0_SDramEn_5, CMOS_DrvX_0_SDramEn_4 => 
        CMOS_DrvX_0_SDramEn_4, CMOS_DrvX_0_SDramEn_3 => 
        CMOS_DrvX_0_SDramEn_3, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[71]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[71]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[70]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[70]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[69]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[69]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[68]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[68]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[67]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[67]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[66]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[66]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[65]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[65]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[64]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[64]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[63]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[63]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[62]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[62]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[61]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[61]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[60]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[60]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[59]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[59]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[58]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[58]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[57]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[57]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[56]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[56]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[55]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[55]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[54]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[54]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[53]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[53]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[52]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[52]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[51]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[51]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[50]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[50]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[49]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[49]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[48]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[48]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[47]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[47]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[46]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[46]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[45]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[45]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[44]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[44]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[43]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[43]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[42]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[42]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[41]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[41]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[40]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[40]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[39]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[39]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[38]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[38]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[37]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[37]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[36]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[36]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[35]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[35]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[34]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[34]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[33]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[33]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[32]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[32]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[31]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[31]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[30]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[30]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[29]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[29]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[28]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[28]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[27]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[27]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[26]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[26]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[25]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[25]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[24]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[24]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[23]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[23]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[22]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[22]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[21]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[21]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[20]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[20]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[19]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[19]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[18]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[18]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[17]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[17]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[16]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[16]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[15]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[15]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[14]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[14]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[13]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[13]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[12]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[12]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[11]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[11]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[10]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[10]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[9]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[9]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[8]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[8]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[7]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[7]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[6]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[6]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[5]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[5]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[4]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[4]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[3]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[3]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[2]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[2]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[1]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[1]\, 
        \Z\\Main_ctl4SD_0_Data2Fifo_[0]\\\ => 
        \Main_ctl4SD_0_Data2Fifo_[0]\, Main_ctl4SD_0_fifo_rst_n
         => Main_ctl4SD_0_fifo_rst_n, FrameMk_0_LVDS_ok => 
        FrameMk_0_LVDS_ok, CMOS_DrvX_0_SDramEn_0 => 
        CMOS_DrvX_0_SDramEn_0, LVDS_enReg => 
        \Sdram_cmd_0.LVDS_enReg\, un6_sdramenreg => 
        \Main_ctl4SD_0.un6_sdramenreg\, CMOS_DrvX_0_AdcEn => 
        CMOS_DrvX_0_AdcEn, N_6 => \Main_ctl4SD_0.N_6\, N_4 => 
        \Main_ctl4SD_0.N_4\, \Z\\My_adder0_0_Sum_[3]\\\ => 
        \My_adder0_0_Sum_[3]\, \Z\\My_adder0_0_Sum_[2]\\\ => 
        \My_adder0_0_Sum_[2]\, \Z\\My_adder0_0_Sum_[1]\\\ => 
        \My_adder0_0_Sum_[1]\, \Z\\My_adder0_0_Sum_[0]\\\ => 
        \My_adder0_0_Sum_[0]\, \Z\\My_adder0_0_Sum_[7]\\\ => 
        \My_adder0_0_Sum_[7]\, \Z\\My_adder0_0_Sum_[6]\\\ => 
        \My_adder0_0_Sum_[6]\, \Z\\My_adder0_0_Sum_[5]\\\ => 
        \My_adder0_0_Sum_[5]\, \Z\\My_adder0_0_Sum_[4]\\\ => 
        \My_adder0_0_Sum_[4]\, \Z\\My_adder0_0_Sum_[11]\\\ => 
        \My_adder0_0_Sum_[11]\, \Z\\My_adder0_0_Sum_[10]\\\ => 
        \My_adder0_0_Sum_[10]\, \Z\\My_adder0_0_Sum_[9]\\\ => 
        \My_adder0_0_Sum_[9]\, \Z\\My_adder0_0_Sum_[8]\\\ => 
        \My_adder0_0_Sum_[8]\, \Z\\My_adder0_0_Sum_[15]\\\ => 
        \My_adder0_0_Sum_[15]\, \Z\\My_adder0_0_Sum_[14]\\\ => 
        \My_adder0_0_Sum_[14]\, \Z\\My_adder0_0_Sum_[13]\\\ => 
        \My_adder0_0_Sum_[13]\, \Z\\My_adder0_0_Sum_[12]\\\ => 
        \My_adder0_0_Sum_[12]\, \Z\\My_adder0_2_Sum_[1]\\\ => 
        \My_adder0_2_Sum_[1]\, \Z\\My_adder0_2_Sum_[0]\\\ => 
        \My_adder0_2_Sum_[0]\, \Z\\My_adder0_1_Sum_[8]\\\ => 
        \My_adder0_1_Sum_[8]\, \Z\\My_adder0_0_Sum_[16]\\\ => 
        \My_adder0_0_Sum_[16]\, \Z\\My_adder0_2_Sum_[3]\\\ => 
        \My_adder0_2_Sum_[3]\, \Z\\My_adder0_2_Sum_[2]\\\ => 
        \My_adder0_2_Sum_[2]\, \Z\\My_adder0_1_Sum_[9]\\\ => 
        \My_adder0_1_Sum_[9]\, \Z\\My_adder0_0_Sum_[17]\\\ => 
        \My_adder0_0_Sum_[17]\, \Z\\My_adder0_2_Sum_[5]\\\ => 
        \My_adder0_2_Sum_[5]\, \Z\\My_adder0_2_Sum_[4]\\\ => 
        \My_adder0_2_Sum_[4]\, \Z\\My_adder0_1_Sum_[10]\\\ => 
        \My_adder0_1_Sum_[10]\, \Z\\My_adder0_1_Sum_[0]\\\ => 
        \My_adder0_1_Sum_[0]\, \Z\\My_adder0_2_Sum_[7]\\\ => 
        \My_adder0_2_Sum_[7]\, \Z\\My_adder0_2_Sum_[6]\\\ => 
        \My_adder0_2_Sum_[6]\, \Z\\My_adder0_1_Sum_[11]\\\ => 
        \My_adder0_1_Sum_[11]\, \Z\\My_adder0_1_Sum_[1]\\\ => 
        \My_adder0_1_Sum_[1]\, \Z\\My_adder0_2_Sum_[9]\\\ => 
        \My_adder0_2_Sum_[9]\, \Z\\My_adder0_2_Sum_[8]\\\ => 
        \My_adder0_2_Sum_[8]\, \Z\\My_adder0_1_Sum_[12]\\\ => 
        \My_adder0_1_Sum_[12]\, \Z\\My_adder0_1_Sum_[2]\\\ => 
        \My_adder0_1_Sum_[2]\, \Z\\My_adder0_2_Sum_[11]\\\ => 
        \My_adder0_2_Sum_[11]\, \Z\\My_adder0_2_Sum_[10]\\\ => 
        \My_adder0_2_Sum_[10]\, \Z\\My_adder0_1_Sum_[13]\\\ => 
        \My_adder0_1_Sum_[13]\, \Z\\My_adder0_1_Sum_[3]\\\ => 
        \My_adder0_1_Sum_[3]\, \Z\\My_adder0_2_Sum_[13]\\\ => 
        \My_adder0_2_Sum_[13]\, \Z\\My_adder0_2_Sum_[12]\\\ => 
        \My_adder0_2_Sum_[12]\, \Z\\My_adder0_1_Sum_[14]\\\ => 
        \My_adder0_1_Sum_[14]\, \Z\\My_adder0_1_Sum_[4]\\\ => 
        \My_adder0_1_Sum_[4]\, \Z\\My_adder0_2_Sum_[15]\\\ => 
        \My_adder0_2_Sum_[15]\, \Z\\My_adder0_2_Sum_[14]\\\ => 
        \My_adder0_2_Sum_[14]\, \Z\\My_adder0_1_Sum_[15]\\\ => 
        \My_adder0_1_Sum_[15]\, \Z\\My_adder0_1_Sum_[5]\\\ => 
        \My_adder0_1_Sum_[5]\, \Z\\My_adder0_2_Sum_[17]\\\ => 
        \My_adder0_2_Sum_[17]\, \Z\\My_adder0_2_Sum_[16]\\\ => 
        \My_adder0_2_Sum_[16]\, \Z\\My_adder0_1_Sum_[16]\\\ => 
        \My_adder0_1_Sum_[16]\, \Z\\My_adder0_1_Sum_[6]\\\ => 
        \My_adder0_1_Sum_[6]\, \Z\\My_adder0_3_Sum_[1]\\\ => 
        \My_adder0_3_Sum_[1]\, \Z\\My_adder0_3_Sum_[0]\\\ => 
        \My_adder0_3_Sum_[0]\, \Z\\My_adder0_1_Sum_[17]\\\ => 
        \My_adder0_1_Sum_[17]\, \Z\\My_adder0_1_Sum_[7]\\\ => 
        \My_adder0_1_Sum_[7]\, \Z\\My_adder0_3_Sum_[5]\\\ => 
        \My_adder0_3_Sum_[5]\, \Z\\My_adder0_3_Sum_[4]\\\ => 
        \My_adder0_3_Sum_[4]\, \Z\\My_adder0_3_Sum_[3]\\\ => 
        \My_adder0_3_Sum_[3]\, \Z\\My_adder0_3_Sum_[2]\\\ => 
        \My_adder0_3_Sum_[2]\, \Z\\My_adder0_3_Sum_[9]\\\ => 
        \My_adder0_3_Sum_[9]\, \Z\\My_adder0_3_Sum_[8]\\\ => 
        \My_adder0_3_Sum_[8]\, \Z\\My_adder0_3_Sum_[7]\\\ => 
        \My_adder0_3_Sum_[7]\, \Z\\My_adder0_3_Sum_[6]\\\ => 
        \My_adder0_3_Sum_[6]\, \Z\\My_adder0_3_Sum_[13]\\\ => 
        \My_adder0_3_Sum_[13]\, \Z\\My_adder0_3_Sum_[12]\\\ => 
        \My_adder0_3_Sum_[12]\, \Z\\My_adder0_3_Sum_[11]\\\ => 
        \My_adder0_3_Sum_[11]\, \Z\\My_adder0_3_Sum_[10]\\\ => 
        \My_adder0_3_Sum_[10]\, \Z\\My_adder0_3_Sum_[17]\\\ => 
        \My_adder0_3_Sum_[17]\, \Z\\My_adder0_3_Sum_[16]\\\ => 
        \My_adder0_3_Sum_[16]\, \Z\\My_adder0_3_Sum_[15]\\\ => 
        \My_adder0_3_Sum_[15]\, \Z\\My_adder0_3_Sum_[14]\\\ => 
        \My_adder0_3_Sum_[14]\, FrameMk_0_LVDS_ok_i => 
        FrameMk_0_LVDS_ok_i, Main_ctl4SD_0_fifo_rst_n_0 => 
        Main_ctl4SD_0_fifo_rst_n_0, Main_ctl4SD_0_fifo_rst_n_1
         => Main_ctl4SD_0_fifo_rst_n_1, 
        Main_ctl4SD_0_fifo_rst_n_2 => Main_ctl4SD_0_fifo_rst_n_2, 
        Main_ctl4SD_0_fifo_rst_n_3 => Main_ctl4SD_0_fifo_rst_n_3, 
        Main_ctl4SD_0_fifo_rst_n_4 => Main_ctl4SD_0_fifo_rst_n_4, 
        Main_ctl4SD_0_fifo_rst_n_5 => Main_ctl4SD_0_fifo_rst_n_5, 
        PLL_Test1_0_SysRst_O => PLL_Test1_0_SysRst_O, 
        PLL_Test1_0_Sys_66M_Clk => PLL_Test1_0_Sys_66M_Clk, 
        Main_ctl4SD_0_fifo_rst_n_6 => Main_ctl4SD_0_fifo_rst_n_6);
    
    \SD_dqm_pad[7]\ : OUTBUF
      port map(D => \SD_dqm_c_c_c_c_c_c_c_c[1]\, PAD => SD_dqm(7));
    
    \SD_dqm_pad[3]\ : OUTBUF
      port map(D => \SD_dqm_c_c_c_c_c_c_c_c[1]\, PAD => SD_dqm(3));
    
    tok_pad : OUTBUF
      port map(D => tok_c, PAD => tok);
    
    \Sd_DQ_pad[34]\ : BIBUF
      port map(PAD => Sd_DQ(34), D => \Fifo_wr_0_Q_[34]\, E => 
        \Sdram_cmd_0.N_264_1\, Y => \Sd_DQ_in[34]\);
    
    \SD_addr_pad[1]\ : OUTBUF
      port map(D => \SD_addr_c[1]\, PAD => SD_addr(1));
    
    spi_load_pad : OUTBUF
      port map(D => spi_load_c, PAD => spi_load);
    
    Pre_co_pad : OUTBUF
      port map(D => Pre_co_c, PAD => Pre_co);
    
    \Sd_DQ_pad[6]\ : BIBUF
      port map(PAD => Sd_DQ(6), D => \Fifo_wr_0_Q_[6]\, E => 
        \Sdram_cmd_0.N_264\, Y => \Sd_DQ_in[6]\);
    
    \Sd_DQ_pad[45]\ : BIBUF
      port map(PAD => Sd_DQ(45), D => \Fifo_wr_0_Q_[45]\, E => 
        \Sdram_cmd_0.N_264_2\, Y => \Sd_DQ_in[45]\);
    
    GND_i_0 : GND
      port map(Y => GND_0);
    
    \Sd_DQ_pad[17]\ : BIBUF
      port map(PAD => Sd_DQ(17), D => \Fifo_wr_0_Q_[17]\, E => 
        \Sdram_cmd_0.N_264_0\, Y => \Sd_DQ_in[17]\);
    
    \SD_addr_pad[12]\ : OUTBUF
      port map(D => \SD_addr_c[12]\, PAD => SD_addr(12));
    
    \Sd_DQ_pad[53]\ : BIBUF
      port map(PAD => Sd_DQ(53), D => \Fifo_wr_0_Q_[53]\, E => 
        \Sdram_cmd_0.N_264_2\, Y => \Sd_DQ_in[53]\);
    
    \SD_addr_pad[10]\ : OUTBUF
      port map(D => \SD_addr_c[10]\, PAD => SD_addr(10));
    
    Fifo_rd_0 : Fifo_rd_1
      port map(\Z\\Fifo_rd_0_Q_[27]\\\ => \Fifo_rd_0_Q_[27]\, 
        \Z\\Fifo_rd_0_Q_[23]\\\ => \Fifo_rd_0_Q_[23]\, 
        \Z\\Fifo_rd_0_Q_[69]\\\ => \Fifo_rd_0_Q_[69]\, 
        \Z\\Fifo_rd_0_Q_[1]\\\ => \Fifo_rd_0_Q_[1]\, 
        \Z\\Fifo_rd_0_Q_[67]\\\ => \Fifo_rd_0_Q_[67]\, 
        \Z\\Fifo_rd_0_Q_[4]\\\ => \Fifo_rd_0_Q_[4]\, 
        \Z\\Fifo_rd_0_Q_[63]\\\ => \Fifo_rd_0_Q_[63]\, 
        \Z\\Fifo_rd_0_Q_[7]\\\ => \Fifo_rd_0_Q_[7]\, 
        \Z\\Fifo_rd_0_Q_[56]\\\ => \Fifo_rd_0_Q_[56]\, 
        \Z\\Fifo_rd_0_Q_[25]\\\ => \Fifo_rd_0_Q_[25]\, 
        \Z\\Fifo_rd_0_Q_[24]\\\ => \Fifo_rd_0_Q_[24]\, 
        \Z\\Fifo_rd_0_Q_[48]\\\ => \Fifo_rd_0_Q_[48]\, 
        \Z\\Fifo_rd_0_Q_[65]\\\ => \Fifo_rd_0_Q_[65]\, 
        \Z\\Fifo_rd_0_Q_[64]\\\ => \Fifo_rd_0_Q_[64]\, 
        \Z\\Fifo_rd_0_Q_[51]\\\ => \Fifo_rd_0_Q_[51]\, 
        \Z\\Fifo_rd_0_Q_[38]\\\ => \Fifo_rd_0_Q_[38]\, 
        \Z\\Fifo_rd_0_Q_[71]\\\ => \Fifo_rd_0_Q_[71]\, 
        \Z\\Fifo_rd_0_Q_[50]\\\ => \Fifo_rd_0_Q_[50]\, 
        \Z\\Fifo_rd_0_Q_[70]\\\ => \Fifo_rd_0_Q_[70]\, 
        \Z\\Fifo_rd_0_Q_[18]\\\ => \Fifo_rd_0_Q_[18]\, 
        \Z\\Fifo_rd_0_Q_[6]\\\ => \Fifo_rd_0_Q_[6]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[71]\\\ => 
        \Sdram_data_0_Sys_dataOut_[71]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[70]\\\ => 
        \Sdram_data_0_Sys_dataOut_[70]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[69]\\\ => 
        \Sdram_data_0_Sys_dataOut_[69]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[68]\\\ => 
        \Sdram_data_0_Sys_dataOut_[68]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[67]\\\ => 
        \Sdram_data_0_Sys_dataOut_[67]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[66]\\\ => 
        \Sdram_data_0_Sys_dataOut_[66]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[65]\\\ => 
        \Sdram_data_0_Sys_dataOut_[65]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[64]\\\ => 
        \Sdram_data_0_Sys_dataOut_[64]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[63]\\\ => 
        \Sdram_data_0_Sys_dataOut_[63]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[62]\\\ => 
        \Sdram_data_0_Sys_dataOut_[62]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[61]\\\ => 
        \Sdram_data_0_Sys_dataOut_[61]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[60]\\\ => 
        \Sdram_data_0_Sys_dataOut_[60]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[59]\\\ => 
        \Sdram_data_0_Sys_dataOut_[59]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[58]\\\ => 
        \Sdram_data_0_Sys_dataOut_[58]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[57]\\\ => 
        \Sdram_data_0_Sys_dataOut_[57]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[56]\\\ => 
        \Sdram_data_0_Sys_dataOut_[56]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[55]\\\ => 
        \Sdram_data_0_Sys_dataOut_[55]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[54]\\\ => 
        \Sdram_data_0_Sys_dataOut_[54]\, \Z\\Fifo_rd_0_Q_[46]\\\
         => \Fifo_rd_0_Q_[46]\, \Z\\Fifo_rd_0_Q_[52]\\\ => 
        \Fifo_rd_0_Q_[52]\, \Z\\Fifo_rd_0_Q_[36]\\\ => 
        \Fifo_rd_0_Q_[36]\, \Z\\Fifo_rd_0_Q_[59]\\\ => 
        \Fifo_rd_0_Q_[59]\, \Z\\Fifo_rd_0_Q_[0]\\\ => 
        \Fifo_rd_0_Q_[0]\, \Z\\Fifo_rd_0_Q_[16]\\\ => 
        \Fifo_rd_0_Q_[16]\, \Z\\Fifo_rd_0_Q_[57]\\\ => 
        \Fifo_rd_0_Q_[57]\, \Z\\Fifo_rd_0_Q_[41]\\\ => 
        \Fifo_rd_0_Q_[41]\, \Z\\Fifo_rd_0_Q_[53]\\\ => 
        \Fifo_rd_0_Q_[53]\, \Z\\Fifo_rd_0_Q_[40]\\\ => 
        \Fifo_rd_0_Q_[40]\, Main_ctl4SD_0_fifo_rd => 
        Main_ctl4SD_0_fifo_rd, \Z\\Fifo_rd_0_Q_[31]\\\ => 
        \Fifo_rd_0_Q_[31]\, \Z\\Fifo_rd_0_Q_[28]\\\ => 
        \Fifo_rd_0_Q_[28]\, \Z\\Fifo_rd_0_Q_[30]\\\ => 
        \Fifo_rd_0_Q_[30]\, \Z\\Fifo_rd_0_Q_[42]\\\ => 
        \Fifo_rd_0_Q_[42]\, \Z\\Fifo_rd_0_Q_[11]\\\ => 
        \Fifo_rd_0_Q_[11]\, \Z\\Fifo_rd_0_Q_[10]\\\ => 
        \Fifo_rd_0_Q_[10]\, \Z\\Fifo_rd_0_Q_[55]\\\ => 
        \Fifo_rd_0_Q_[55]\, \Z\\Fifo_rd_0_Q_[68]\\\ => 
        \Fifo_rd_0_Q_[68]\, \Z\\Fifo_rd_0_Q_[54]\\\ => 
        \Fifo_rd_0_Q_[54]\, \Z\\Fifo_rd_0_Q_[49]\\\ => 
        \Fifo_rd_0_Q_[49]\, \Z\\Fifo_rd_0_Q_[9]\\\ => 
        \Fifo_rd_0_Q_[9]\, \Z\\Fifo_rd_0_Q_[5]\\\ => 
        \Fifo_rd_0_Q_[5]\, Fifo_rd_0_AFULL => Fifo_rd_0_AFULL, 
        \Z\\Fifo_rd_0_Q_[32]\\\ => \Fifo_rd_0_Q_[32]\, 
        \Z\\Fifo_rd_0_Q_[47]\\\ => \Fifo_rd_0_Q_[47]\, 
        \Z\\Fifo_rd_0_Q_[43]\\\ => \Fifo_rd_0_Q_[43]\, 
        \Z\\Fifo_rd_0_Q_[12]\\\ => \Fifo_rd_0_Q_[12]\, 
        Sdram_cmd_0_RFifo_we => Sdram_cmd_0_RFifo_we, 
        \Z\\Fifo_rd_0_Q_[26]\\\ => \Fifo_rd_0_Q_[26]\, 
        \Z\\Fifo_rd_0_Q_[39]\\\ => \Fifo_rd_0_Q_[39]\, 
        \Z\\Fifo_rd_0_Q_[19]\\\ => \Fifo_rd_0_Q_[19]\, 
        \Z\\Fifo_rd_0_Q_[37]\\\ => \Fifo_rd_0_Q_[37]\, 
        \Z\\Fifo_rd_0_Q_[3]\\\ => \Fifo_rd_0_Q_[3]\, 
        \Z\\Fifo_rd_0_Q_[33]\\\ => \Fifo_rd_0_Q_[33]\, 
        \Z\\Fifo_rd_0_Q_[66]\\\ => \Fifo_rd_0_Q_[66]\, 
        \Z\\Fifo_rd_0_Q_[17]\\\ => \Fifo_rd_0_Q_[17]\, 
        \Z\\Fifo_rd_0_Q_[13]\\\ => \Fifo_rd_0_Q_[13]\, 
        \Z\\Fifo_rd_0_Q_[45]\\\ => \Fifo_rd_0_Q_[45]\, 
        \Z\\Fifo_rd_0_Q_[44]\\\ => \Fifo_rd_0_Q_[44]\, 
        \Z\\Fifo_rd_0_Q_[21]\\\ => \Fifo_rd_0_Q_[21]\, 
        \Z\\Fifo_rd_0_Q_[2]\\\ => \Fifo_rd_0_Q_[2]\, 
        \Z\\Fifo_rd_0_Q_[20]\\\ => \Fifo_rd_0_Q_[20]\, 
        \Z\\Fifo_rd_0_Q_[61]\\\ => \Fifo_rd_0_Q_[61]\, 
        \Z\\Fifo_rd_0_Q_[35]\\\ => \Fifo_rd_0_Q_[35]\, 
        \Z\\Fifo_rd_0_Q_[34]\\\ => \Fifo_rd_0_Q_[34]\, 
        \Z\\Fifo_rd_0_Q_[60]\\\ => \Fifo_rd_0_Q_[60]\, 
        \Z\\Fifo_rd_0_Q_[15]\\\ => \Fifo_rd_0_Q_[15]\, 
        \Z\\Fifo_rd_0_Q_[14]\\\ => \Fifo_rd_0_Q_[14]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[35]\\\ => 
        \Sdram_data_0_Sys_dataOut_[35]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[34]\\\ => 
        \Sdram_data_0_Sys_dataOut_[34]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[33]\\\ => 
        \Sdram_data_0_Sys_dataOut_[33]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[32]\\\ => 
        \Sdram_data_0_Sys_dataOut_[32]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[31]\\\ => 
        \Sdram_data_0_Sys_dataOut_[31]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[30]\\\ => 
        \Sdram_data_0_Sys_dataOut_[30]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[29]\\\ => 
        \Sdram_data_0_Sys_dataOut_[29]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[28]\\\ => 
        \Sdram_data_0_Sys_dataOut_[28]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[27]\\\ => 
        \Sdram_data_0_Sys_dataOut_[27]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[26]\\\ => 
        \Sdram_data_0_Sys_dataOut_[26]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[25]\\\ => 
        \Sdram_data_0_Sys_dataOut_[25]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[24]\\\ => 
        \Sdram_data_0_Sys_dataOut_[24]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[23]\\\ => 
        \Sdram_data_0_Sys_dataOut_[23]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[22]\\\ => 
        \Sdram_data_0_Sys_dataOut_[22]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[21]\\\ => 
        \Sdram_data_0_Sys_dataOut_[21]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[20]\\\ => 
        \Sdram_data_0_Sys_dataOut_[20]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[19]\\\ => 
        \Sdram_data_0_Sys_dataOut_[19]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[18]\\\ => 
        \Sdram_data_0_Sys_dataOut_[18]\, 
        Main_ctl4SD_0_fifo_rst_n_0 => Main_ctl4SD_0_fifo_rst_n_0, 
        \Z\\Fifo_rd_0_Q_[22]\\\ => \Fifo_rd_0_Q_[22]\, 
        \Z\\Fifo_rd_0_Q_[8]\\\ => \Fifo_rd_0_Q_[8]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[53]\\\ => 
        \Sdram_data_0_Sys_dataOut_[53]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[52]\\\ => 
        \Sdram_data_0_Sys_dataOut_[52]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[51]\\\ => 
        \Sdram_data_0_Sys_dataOut_[51]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[50]\\\ => 
        \Sdram_data_0_Sys_dataOut_[50]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[49]\\\ => 
        \Sdram_data_0_Sys_dataOut_[49]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[48]\\\ => 
        \Sdram_data_0_Sys_dataOut_[48]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[47]\\\ => 
        \Sdram_data_0_Sys_dataOut_[47]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[46]\\\ => 
        \Sdram_data_0_Sys_dataOut_[46]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[45]\\\ => 
        \Sdram_data_0_Sys_dataOut_[45]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[44]\\\ => 
        \Sdram_data_0_Sys_dataOut_[44]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[43]\\\ => 
        \Sdram_data_0_Sys_dataOut_[43]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[42]\\\ => 
        \Sdram_data_0_Sys_dataOut_[42]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[41]\\\ => 
        \Sdram_data_0_Sys_dataOut_[41]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[40]\\\ => 
        \Sdram_data_0_Sys_dataOut_[40]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[39]\\\ => 
        \Sdram_data_0_Sys_dataOut_[39]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[38]\\\ => 
        \Sdram_data_0_Sys_dataOut_[38]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[37]\\\ => 
        \Sdram_data_0_Sys_dataOut_[37]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[36]\\\ => 
        \Sdram_data_0_Sys_dataOut_[36]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[17]\\\ => 
        \Sdram_data_0_Sys_dataOut_[17]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[16]\\\ => 
        \Sdram_data_0_Sys_dataOut_[16]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[15]\\\ => 
        \Sdram_data_0_Sys_dataOut_[15]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[14]\\\ => 
        \Sdram_data_0_Sys_dataOut_[14]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[13]\\\ => 
        \Sdram_data_0_Sys_dataOut_[13]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[12]\\\ => 
        \Sdram_data_0_Sys_dataOut_[12]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[11]\\\ => 
        \Sdram_data_0_Sys_dataOut_[11]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[10]\\\ => 
        \Sdram_data_0_Sys_dataOut_[10]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[9]\\\ => 
        \Sdram_data_0_Sys_dataOut_[9]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[8]\\\ => 
        \Sdram_data_0_Sys_dataOut_[8]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[7]\\\ => 
        \Sdram_data_0_Sys_dataOut_[7]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[6]\\\ => 
        \Sdram_data_0_Sys_dataOut_[6]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[5]\\\ => 
        \Sdram_data_0_Sys_dataOut_[5]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[4]\\\ => 
        \Sdram_data_0_Sys_dataOut_[4]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[3]\\\ => 
        \Sdram_data_0_Sys_dataOut_[3]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[2]\\\ => 
        \Sdram_data_0_Sys_dataOut_[2]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[1]\\\ => 
        \Sdram_data_0_Sys_dataOut_[1]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[0]\\\ => 
        \Sdram_data_0_Sys_dataOut_[0]\, Fifo_rd_1_VCC => \VCC\, 
        Main_ctl4SD_0_fifo_rst_n_3 => Main_ctl4SD_0_fifo_rst_n_3, 
        \Z\\Fifo_rd_0_Q_[62]\\\ => \Fifo_rd_0_Q_[62]\, 
        Main_ctl4SD_0_fifo_rst_n_1 => Main_ctl4SD_0_fifo_rst_n_1, 
        \Z\\Fifo_rd_0_Q_[29]\\\ => \Fifo_rd_0_Q_[29]\, 
        Main_ctl4SD_0_fifo_rst_n_2 => Main_ctl4SD_0_fifo_rst_n_2, 
        PLL_Test1_0_Sys_66M_Clk => PLL_Test1_0_Sys_66M_Clk, 
        \Z\\Fifo_rd_0_Q_[58]\\\ => \Fifo_rd_0_Q_[58]\, 
        Fifo_rd_1_GND => \GND\);
    
    \Sd_DQ_pad[27]\ : BIBUF
      port map(PAD => Sd_DQ(27), D => \Fifo_wr_0_Q_[27]\, E => 
        \Sdram_cmd_0.N_264_1\, Y => \Sd_DQ_in[27]\);
    
    spi_data_pad : OUTBUF
      port map(D => spi_data_c, PAD => spi_data);
    
    \SD_addr_pad[6]\ : OUTBUF
      port map(D => \SD_addr_c[6]\, PAD => SD_addr(6));
    
    \Sd_DQ_pad[44]\ : BIBUF
      port map(PAD => Sd_DQ(44), D => \Fifo_wr_0_Q_[44]\, E => 
        \Sdram_cmd_0.N_264_2\, Y => \Sd_DQ_in[44]\);
    
    Prebus2_pad : OUTBUF
      port map(D => \GND\, PAD => Prebus2);
    
    \SD_dqm_pad[0]\ : OUTBUF
      port map(D => \SD_dqm_c_c_c_c_c_c_c_c[1]\, PAD => SD_dqm(0));
    
    \SD_dqm_pad[6]\ : OUTBUF
      port map(D => \SD_dqm_c_c_c_c_c_c_c_c[1]\, PAD => SD_dqm(6));
    
    \SD_addr_pad[5]\ : OUTBUF
      port map(D => \SD_addr_c[5]\, PAD => SD_addr(5));
    
    Sdram_data_0 : Sdram_data
      port map(Sd_DQ_in(71) => \Sd_DQ_in[71]\, Sd_DQ_in(70) => 
        \Sd_DQ_in[70]\, Sd_DQ_in(69) => \Sd_DQ_in[69]\, 
        Sd_DQ_in(68) => \Sd_DQ_in[68]\, Sd_DQ_in(67) => 
        \Sd_DQ_in[67]\, Sd_DQ_in(66) => \Sd_DQ_in[66]\, 
        Sd_DQ_in(65) => \Sd_DQ_in[65]\, Sd_DQ_in(64) => 
        \Sd_DQ_in[64]\, Sd_DQ_in(63) => \Sd_DQ_in[63]\, 
        Sd_DQ_in(62) => \Sd_DQ_in[62]\, Sd_DQ_in(61) => 
        \Sd_DQ_in[61]\, Sd_DQ_in(60) => \Sd_DQ_in[60]\, 
        Sd_DQ_in(59) => \Sd_DQ_in[59]\, Sd_DQ_in(58) => 
        \Sd_DQ_in[58]\, Sd_DQ_in(57) => \Sd_DQ_in[57]\, 
        Sd_DQ_in(56) => \Sd_DQ_in[56]\, Sd_DQ_in(55) => 
        \Sd_DQ_in[55]\, Sd_DQ_in(54) => \Sd_DQ_in[54]\, 
        Sd_DQ_in(53) => \Sd_DQ_in[53]\, Sd_DQ_in(52) => 
        \Sd_DQ_in[52]\, Sd_DQ_in(51) => \Sd_DQ_in[51]\, 
        Sd_DQ_in(50) => \Sd_DQ_in[50]\, Sd_DQ_in(49) => 
        \Sd_DQ_in[49]\, Sd_DQ_in(48) => \Sd_DQ_in[48]\, 
        Sd_DQ_in(47) => \Sd_DQ_in[47]\, Sd_DQ_in(46) => 
        \Sd_DQ_in[46]\, Sd_DQ_in(45) => \Sd_DQ_in[45]\, 
        Sd_DQ_in(44) => \Sd_DQ_in[44]\, Sd_DQ_in(43) => 
        \Sd_DQ_in[43]\, Sd_DQ_in(42) => \Sd_DQ_in[42]\, 
        Sd_DQ_in(41) => \Sd_DQ_in[41]\, Sd_DQ_in(40) => 
        \Sd_DQ_in[40]\, Sd_DQ_in(39) => \Sd_DQ_in[39]\, 
        Sd_DQ_in(38) => \Sd_DQ_in[38]\, Sd_DQ_in(37) => 
        \Sd_DQ_in[37]\, Sd_DQ_in(36) => \Sd_DQ_in[36]\, 
        Sd_DQ_in(35) => \Sd_DQ_in[35]\, Sd_DQ_in(34) => 
        \Sd_DQ_in[34]\, Sd_DQ_in(33) => \Sd_DQ_in[33]\, 
        Sd_DQ_in(32) => \Sd_DQ_in[32]\, Sd_DQ_in(31) => 
        \Sd_DQ_in[31]\, Sd_DQ_in(30) => \Sd_DQ_in[30]\, 
        Sd_DQ_in(29) => \Sd_DQ_in[29]\, Sd_DQ_in(28) => 
        \Sd_DQ_in[28]\, Sd_DQ_in(27) => \Sd_DQ_in[27]\, 
        Sd_DQ_in(26) => \Sd_DQ_in[26]\, Sd_DQ_in(25) => 
        \Sd_DQ_in[25]\, Sd_DQ_in(24) => \Sd_DQ_in[24]\, 
        Sd_DQ_in(23) => \Sd_DQ_in[23]\, Sd_DQ_in(22) => 
        \Sd_DQ_in[22]\, Sd_DQ_in(21) => \Sd_DQ_in[21]\, 
        Sd_DQ_in(20) => \Sd_DQ_in[20]\, Sd_DQ_in(19) => 
        \Sd_DQ_in[19]\, Sd_DQ_in(18) => \Sd_DQ_in[18]\, 
        Sd_DQ_in(17) => \Sd_DQ_in[17]\, Sd_DQ_in(16) => 
        \Sd_DQ_in[16]\, Sd_DQ_in(15) => \Sd_DQ_in[15]\, 
        Sd_DQ_in(14) => \Sd_DQ_in[14]\, Sd_DQ_in(13) => 
        \Sd_DQ_in[13]\, Sd_DQ_in(12) => \Sd_DQ_in[12]\, 
        Sd_DQ_in(11) => \Sd_DQ_in[11]\, Sd_DQ_in(10) => 
        \Sd_DQ_in[10]\, Sd_DQ_in(9) => \Sd_DQ_in[9]\, Sd_DQ_in(8)
         => \Sd_DQ_in[8]\, Sd_DQ_in(7) => \Sd_DQ_in[7]\, 
        Sd_DQ_in(6) => \Sd_DQ_in[6]\, Sd_DQ_in(5) => 
        \Sd_DQ_in[5]\, Sd_DQ_in(4) => \Sd_DQ_in[4]\, Sd_DQ_in(3)
         => \Sd_DQ_in[3]\, Sd_DQ_in(2) => \Sd_DQ_in[2]\, 
        Sd_DQ_in(1) => \Sd_DQ_in[1]\, Sd_DQ_in(0) => 
        \Sd_DQ_in[0]\, \Z\\Sdram_data_0_Sys_dataOut_[71]\\\ => 
        \Sdram_data_0_Sys_dataOut_[71]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[70]\\\ => 
        \Sdram_data_0_Sys_dataOut_[70]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[69]\\\ => 
        \Sdram_data_0_Sys_dataOut_[69]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[68]\\\ => 
        \Sdram_data_0_Sys_dataOut_[68]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[67]\\\ => 
        \Sdram_data_0_Sys_dataOut_[67]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[66]\\\ => 
        \Sdram_data_0_Sys_dataOut_[66]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[65]\\\ => 
        \Sdram_data_0_Sys_dataOut_[65]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[64]\\\ => 
        \Sdram_data_0_Sys_dataOut_[64]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[63]\\\ => 
        \Sdram_data_0_Sys_dataOut_[63]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[62]\\\ => 
        \Sdram_data_0_Sys_dataOut_[62]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[61]\\\ => 
        \Sdram_data_0_Sys_dataOut_[61]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[60]\\\ => 
        \Sdram_data_0_Sys_dataOut_[60]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[59]\\\ => 
        \Sdram_data_0_Sys_dataOut_[59]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[58]\\\ => 
        \Sdram_data_0_Sys_dataOut_[58]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[57]\\\ => 
        \Sdram_data_0_Sys_dataOut_[57]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[56]\\\ => 
        \Sdram_data_0_Sys_dataOut_[56]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[55]\\\ => 
        \Sdram_data_0_Sys_dataOut_[55]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[54]\\\ => 
        \Sdram_data_0_Sys_dataOut_[54]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[53]\\\ => 
        \Sdram_data_0_Sys_dataOut_[53]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[52]\\\ => 
        \Sdram_data_0_Sys_dataOut_[52]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[51]\\\ => 
        \Sdram_data_0_Sys_dataOut_[51]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[50]\\\ => 
        \Sdram_data_0_Sys_dataOut_[50]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[49]\\\ => 
        \Sdram_data_0_Sys_dataOut_[49]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[48]\\\ => 
        \Sdram_data_0_Sys_dataOut_[48]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[47]\\\ => 
        \Sdram_data_0_Sys_dataOut_[47]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[46]\\\ => 
        \Sdram_data_0_Sys_dataOut_[46]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[45]\\\ => 
        \Sdram_data_0_Sys_dataOut_[45]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[44]\\\ => 
        \Sdram_data_0_Sys_dataOut_[44]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[43]\\\ => 
        \Sdram_data_0_Sys_dataOut_[43]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[42]\\\ => 
        \Sdram_data_0_Sys_dataOut_[42]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[41]\\\ => 
        \Sdram_data_0_Sys_dataOut_[41]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[40]\\\ => 
        \Sdram_data_0_Sys_dataOut_[40]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[39]\\\ => 
        \Sdram_data_0_Sys_dataOut_[39]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[38]\\\ => 
        \Sdram_data_0_Sys_dataOut_[38]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[37]\\\ => 
        \Sdram_data_0_Sys_dataOut_[37]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[36]\\\ => 
        \Sdram_data_0_Sys_dataOut_[36]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[35]\\\ => 
        \Sdram_data_0_Sys_dataOut_[35]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[34]\\\ => 
        \Sdram_data_0_Sys_dataOut_[34]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[33]\\\ => 
        \Sdram_data_0_Sys_dataOut_[33]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[32]\\\ => 
        \Sdram_data_0_Sys_dataOut_[32]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[31]\\\ => 
        \Sdram_data_0_Sys_dataOut_[31]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[30]\\\ => 
        \Sdram_data_0_Sys_dataOut_[30]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[29]\\\ => 
        \Sdram_data_0_Sys_dataOut_[29]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[28]\\\ => 
        \Sdram_data_0_Sys_dataOut_[28]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[27]\\\ => 
        \Sdram_data_0_Sys_dataOut_[27]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[26]\\\ => 
        \Sdram_data_0_Sys_dataOut_[26]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[25]\\\ => 
        \Sdram_data_0_Sys_dataOut_[25]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[24]\\\ => 
        \Sdram_data_0_Sys_dataOut_[24]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[23]\\\ => 
        \Sdram_data_0_Sys_dataOut_[23]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[22]\\\ => 
        \Sdram_data_0_Sys_dataOut_[22]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[21]\\\ => 
        \Sdram_data_0_Sys_dataOut_[21]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[20]\\\ => 
        \Sdram_data_0_Sys_dataOut_[20]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[19]\\\ => 
        \Sdram_data_0_Sys_dataOut_[19]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[18]\\\ => 
        \Sdram_data_0_Sys_dataOut_[18]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[17]\\\ => 
        \Sdram_data_0_Sys_dataOut_[17]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[16]\\\ => 
        \Sdram_data_0_Sys_dataOut_[16]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[15]\\\ => 
        \Sdram_data_0_Sys_dataOut_[15]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[14]\\\ => 
        \Sdram_data_0_Sys_dataOut_[14]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[13]\\\ => 
        \Sdram_data_0_Sys_dataOut_[13]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[12]\\\ => 
        \Sdram_data_0_Sys_dataOut_[12]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[11]\\\ => 
        \Sdram_data_0_Sys_dataOut_[11]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[10]\\\ => 
        \Sdram_data_0_Sys_dataOut_[10]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[9]\\\ => 
        \Sdram_data_0_Sys_dataOut_[9]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[8]\\\ => 
        \Sdram_data_0_Sys_dataOut_[8]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[7]\\\ => 
        \Sdram_data_0_Sys_dataOut_[7]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[6]\\\ => 
        \Sdram_data_0_Sys_dataOut_[6]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[5]\\\ => 
        \Sdram_data_0_Sys_dataOut_[5]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[4]\\\ => 
        \Sdram_data_0_Sys_dataOut_[4]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[3]\\\ => 
        \Sdram_data_0_Sys_dataOut_[3]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[2]\\\ => 
        \Sdram_data_0_Sys_dataOut_[2]\, 
        \Z\\Sdram_data_0_Sys_dataOut_[1]\\\ => 
        \Sdram_data_0_Sys_dataOut_[1]\, PLL_Test1_0_SysRst_O => 
        PLL_Test1_0_SysRst_O, PLL_Test1_0_Sys_66M_Clk => 
        PLL_Test1_0_Sys_66M_Clk, 
        \Z\\Sdram_data_0_Sys_dataOut_[0]\\\ => 
        \Sdram_data_0_Sys_dataOut_[0]\, 
        \Z\\SDram_rd_0_rd_state_[1]\\\ => 
        \SDram_rd_0_rd_state_[1]\, \Z\\SDram_rd_0_rd_state_[2]\\\
         => \SDram_rd_0_rd_state_[2]\, 
        \Z\\SDram_rd_0_rd_state_[0]\\\ => 
        \SDram_rd_0_rd_state_[0]\);
    
    adc_muxtmp_test_0 : adc_muxtmp_test
      port map(PLL_Test1_0_SysRst_O => PLL_Test1_0_SysRst_O, 
        PLL_Test1_0_Sys_66M_Clk => PLL_Test1_0_Sys_66M_Clk, 
        CMOS_DrvX_0_AdcEn => CMOS_DrvX_0_AdcEn, 
        \Z\\adc_muxtmp_test_0_DataOut41to28_[29]\\\ => 
        \adc_muxtmp_test_0_DataOut41to28_[29]\, 
        \Z\\adc_muxtmp_test_0_DataOut27to14_[14]\\\ => 
        \adc_muxtmp_test_0_DataOut27to14_[14]\, 
        \Z\\adc_muxtmp_test_0_DataOut55to42_[43]\\\ => 
        \adc_muxtmp_test_0_DataOut55to42_[43]\);
    
    \Sd_DQ_pad[55]\ : BIBUF
      port map(PAD => Sd_DQ(55), D => \Fifo_wr_0_Q_[55]\, E => 
        \Sdram_cmd_0.N_264_2\, Y => \Sd_DQ_in[55]\);
    
    reset_ds_pad : OUTBUF
      port map(D => \GND\, PAD => reset_ds);
    
    \Sd_DQ_pad[9]\ : BIBUF
      port map(PAD => Sd_DQ(9), D => \Fifo_wr_0_Q_[9]\, E => 
        \Sdram_cmd_0.N_264\, Y => \Sd_DQ_in[9]\);
    
    \Sd_DQ_pad[67]\ : BIBUF
      port map(PAD => Sd_DQ(67), D => \Fifo_wr_0_Q_[67]\, E => 
        \Sdram_cmd_0.N_264\, Y => \Sd_DQ_in[67]\);
    
    PLL_Test1_0 : PLL_Test1
      port map(PLL_Test1_0_ADC_66M_Clk => PLL_Test1_0_ADC_66M_Clk, 
        PLL_Test1_0_Sdram_clk => PLL_Test1_0_Sdram_clk, 
        ExterCLk_c => ExterCLk_c, PLL_Test1_GND => \GND\, 
        PLL_Test1_0_SysRst_O => PLL_Test1_0_SysRst_O, 
        PLL_Test1_VCC => \VCC\, PLL_Test1_0_Sys_66M_Clk => 
        PLL_Test1_0_Sys_66M_Clk);
    
    \Sd_DQ_pad[12]\ : BIBUF
      port map(PAD => Sd_DQ(12), D => \Fifo_wr_0_Q_[12]\, E => 
        \Sdram_cmd_0.N_264_0\, Y => \Sd_DQ_in[12]\);
    
    \SD_Clk_pad[0]\ : OUTBUF
      port map(D => \SD_Clk_c_c[1]\, PAD => SD_Clk(0));
    
    \SD_addr_pad[9]\ : OUTBUF
      port map(D => \SD_addr_c[9]\, PAD => SD_addr(9));
    
    \Sd_DQ_pad[54]\ : BIBUF
      port map(PAD => Sd_DQ(54), D => \Fifo_wr_0_Q_[54]\, E => 
        \Sdram_cmd_0.N_264_2\, Y => \Sd_DQ_in[54]\);
    
    \Sd_DQ_pad[8]\ : BIBUF
      port map(PAD => Sd_DQ(8), D => \Fifo_wr_0_Q_[8]\, E => 
        \Sdram_cmd_0.N_264\, Y => \Sd_DQ_in[8]\);
    
    \Sd_DQ_pad[22]\ : BIBUF
      port map(PAD => Sd_DQ(22), D => \Fifo_wr_0_Q_[22]\, E => 
        \Sdram_cmd_0.N_264_0\, Y => \Sd_DQ_in[22]\);
    
    \Sd_DQ_pad[19]\ : BIBUF
      port map(PAD => Sd_DQ(19), D => \Fifo_wr_0_Q_[19]\, E => 
        \Sdram_cmd_0.N_264_0\, Y => \Sd_DQ_in[19]\);
    
    \Sd_DQ_pad[16]\ : BIBUF
      port map(PAD => Sd_DQ(16), D => \Fifo_wr_0_Q_[16]\, E => 
        \Sdram_cmd_0.N_264_0\, Y => \Sd_DQ_in[16]\);
    
    Sdram_ctl_v2_0 : Sdram_ctl_v2
      port map(SD_cke_c_c(0) => \SD_cke_c_c[0]\, pr_state_ns_3
         => \Sdram_ctl_v2_0.pr_state_ns[8]\, 
        Sdram_ini_0_Sd_iniOK_i => Sdram_ini_0_Sd_iniOK_i, 
        Sdram_ctl_v2_0_SD_iniEn => Sdram_ctl_v2_0_SD_iniEn, 
        Sdram_ctl_v2_0_SD_RefEn => Sdram_ctl_v2_0_SD_RefEn, 
        Sdram_ctl_v2_0_SD_rdEN_noact => 
        Sdram_ctl_v2_0_SD_rdEN_noact, PLL_Test1_0_SysRst_O => 
        PLL_Test1_0_SysRst_O, PLL_Test1_0_Sys_66M_Clk => 
        PLL_Test1_0_Sys_66M_Clk, Sdram_ctl_v2_0_SD_pdEN => 
        Sdram_ctl_v2_0_SD_pdEN, Fifo_wr_0_AFULL => 
        Fifo_wr_0_AFULL, SDRAM_wr_0_SD_WrOK => SDRAM_wr_0_SD_WrOK, 
        ref_ok_2 => \SDRAM_Ref_0.ref_ok_2\, ref_ok_1 => 
        \SDRAM_Ref_0.ref_ok_1\, CMOS_DrvX_0_LVDSen_2 => 
        CMOS_DrvX_0_LVDSen_2, CMOS_DrvX_0_SDramEn_0 => 
        CMOS_DrvX_0_SDramEn_0, Sdram_ini_0_Sd_iniOK => 
        Sdram_ini_0_Sd_iniOK, Fifo_rd_0_AFULL => Fifo_rd_0_AFULL, 
        CMOS_DrvX_0_LVDSen_1 => CMOS_DrvX_0_LVDSen_1, 
        SDram_rd_0_SD_RdOK => SDram_rd_0_SD_RdOK, 
        Sdram_ctl_v2_0_SD_rdEn => Sdram_ctl_v2_0_SD_rdEn, 
        Sdram_ctl_v2_0_SD_rdEn_i => Sdram_ctl_v2_0_SD_rdEn_i, 
        Sdram_ctl_v2_0_SD_wrEn => Sdram_ctl_v2_0_SD_wrEn, 
        Sdram_ctl_v2_0_SD_wrEn_i => Sdram_ctl_v2_0_SD_wrEn_i);
    
    \Sd_DQ_pad[37]\ : BIBUF
      port map(PAD => Sd_DQ(37), D => \Fifo_wr_0_Q_[37]\, E => 
        \Sdram_cmd_0.N_264_1\, Y => \Sd_DQ_in[37]\);
    
    \SD_addr_pad[11]\ : OUTBUF
      port map(D => \SD_addr_c[11]\, PAD => SD_addr(11));
    
    \Sd_DQ_pad[29]\ : BIBUF
      port map(PAD => Sd_DQ(29), D => \Fifo_wr_0_Q_[29]\, E => 
        \Sdram_cmd_0.N_264_1\, Y => \Sd_DQ_in[29]\);
    
    \Sd_DQ_pad[26]\ : BIBUF
      port map(PAD => Sd_DQ(26), D => \Fifo_wr_0_Q_[26]\, E => 
        \Sdram_cmd_0.N_264_1\, Y => \Sd_DQ_in[26]\);
    
    \Sd_DQ_pad[0]\ : BIBUF
      port map(PAD => Sd_DQ(0), D => \Fifo_wr_0_Q_[0]\, E => 
        \Sdram_cmd_0.N_264_0\, Y => \Sd_DQ_in[0]\);
    
    \Sd_DQ_pad[10]\ : BIBUF
      port map(PAD => Sd_DQ(10), D => \Fifo_wr_0_Q_[10]\, E => 
        \Sdram_cmd_0.N_264_0\, Y => \Sd_DQ_in[10]\);
    
    \My_adder0_1\ : My_adder0_2
      port map(intData2acc_RNI2KS7(28) => 
        \intData2acc_RNI2KS7[28]\, intData2acc_RNI1KS7(27) => 
        \intData2acc_RNI1KS7[27]\, intData2acc_RNI6JV9(33) => 
        \intData2acc_RNI6JV9[33]\, intData2acc_RNI2BV9(18) => 
        \intData2acc_RNI2BV9[18]\, intData2acc_RNI3BV9(19) => 
        \intData2acc_RNI3BV9[19]\, intData2acc_RNIBN36(22) => 
        \intData2acc_RNIBN36[22]\, intData2acc_RNI3JV9(30) => 
        \intData2acc_RNI3JV9[30]\, intData2acc_RNI5JV9(32) => 
        \intData2acc_RNI5JV9[32]\, intData2acc_RNITEV9(20) => 
        \intData2acc_RNITEV9[20]\, intData2acc_RNIAN36(21) => 
        \intData2acc_RNIAN36[21]\, intData2acc_RNI4JV9(31) => 
        \intData2acc_RNI4JV9[31]\, intData2acc_RNIDN36(24) => 
        \intData2acc_RNIDN36[24]\, intData2acc_RNIEN36(25) => 
        \intData2acc_RNIEN36[25]\, intData2acc_RNI9FV9(29) => 
        \intData2acc_RNI9FV9[29]\, intData2acc_RNI8JV9(35) => 
        \intData2acc_RNI8JV9[35]\, intData2acc_RNITJS7(23) => 
        \intData2acc_RNITJS7[23]\, intData2acc_RNI0KS7(26) => 
        \intData2acc_RNI0KS7[26]\, intData2acc_RNI7JV9(34) => 
        \intData2acc_RNI7JV9[34]\, \Z\\My_adder0_1_Sum_[15]\\\
         => \My_adder0_1_Sum_[15]\, \Z\\My_adder0_1_Sum_[12]\\\
         => \My_adder0_1_Sum_[12]\, \Z\\My_adder0_1_Sum_[6]\\\
         => \My_adder0_1_Sum_[6]\, \Z\\My_adder0_1_Sum_[10]\\\
         => \My_adder0_1_Sum_[10]\, \Z\\My_adder0_1_Sum_[9]\\\
         => \My_adder0_1_Sum_[9]\, \Z\\My_adder0_1_Sum_[7]\\\ => 
        \My_adder0_1_Sum_[7]\, \Z\\My_adder0_1_Sum_[11]\\\ => 
        \My_adder0_1_Sum_[11]\, \Z\\My_adder0_1_Sum_[1]\\\ => 
        \My_adder0_1_Sum_[1]\, \Z\\My_adder0_1_Sum_[3]\\\ => 
        \My_adder0_1_Sum_[3]\, \Z\\My_adder0_1_Sum_[13]\\\ => 
        \My_adder0_1_Sum_[13]\, 
        \Z\\adc_muxtmp_test_0_DataOut27to14_[14]\\\ => 
        \adc_muxtmp_test_0_DataOut27to14_[14]\, 
        \Z\\My_adder0_1_Sum_[0]\\\ => \My_adder0_1_Sum_[0]\, 
        \Z\\My_adder0_1_Sum_[8]\\\ => \My_adder0_1_Sum_[8]\, 
        \Z\\My_adder0_1_Sum_[14]\\\ => \My_adder0_1_Sum_[14]\, 
        \Z\\My_adder0_1_Sum_[2]\\\ => \My_adder0_1_Sum_[2]\, 
        \Z\\My_adder0_1_Sum_[4]\\\ => \My_adder0_1_Sum_[4]\, 
        \Z\\My_adder0_1_Sum_[5]\\\ => \My_adder0_1_Sum_[5]\, 
        \Z\\My_adder0_1_Sum_[17]\\\ => \My_adder0_1_Sum_[17]\, 
        My_adder0_2_GND => \GND\, \Z\\My_adder0_1_Sum_[16]\\\ => 
        \My_adder0_1_Sum_[16]\);
    
    Clock_Y_pad : OUTBUF
      port map(D => Clock_Y_c, PAD => Clock_Y);
    
    \Sd_DQ_pad[20]\ : BIBUF
      port map(PAD => Sd_DQ(20), D => \Fifo_wr_0_Q_[20]\, E => 
        \Sdram_cmd_0.N_264_0\, Y => \Sd_DQ_in[20]\);
    
    \Sd_DQ_pad[7]\ : BIBUF
      port map(PAD => Sd_DQ(7), D => \Fifo_wr_0_Q_[7]\, E => 
        \Sdram_cmd_0.N_264\, Y => \Sd_DQ_in[7]\);
    
    VoltAvg_pad : OUTBUF
      port map(D => \GND\, PAD => VoltAvg);
    
    \Sd_DQ_pad[18]\ : BIBUF
      port map(PAD => Sd_DQ(18), D => \Fifo_wr_0_Q_[18]\, E => 
        \Sdram_cmd_0.N_264_0\, Y => \Sd_DQ_in[18]\);
    

end DEF_ARCH; 
